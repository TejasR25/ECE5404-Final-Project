//`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.05.2024 04:35:38
// Design Name: 
// Module Name: pca_score
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module min_pca_score
#(
    parameter MIN_PC_NUM = 5) 
    
    (
//********************************************************* USING 64 BIT BINARY *********************************************************************
//---------------------------------------------- CLOCK INSERTED ----------------------------------------------------------
 //   input wire clk, reset,
//    input wire [FP_SIZE-1:0] min_eigen_values [0:MIN_PC_NUM-1],
//    input wire [FP_SIZE-1:0] min_principal_comps [0:MIN_PC_NUM-1],
//    output wire [FP_SIZE-1:0] min_pc_score
//------------------------------------------------------------------------------------------------------------------------
//---------------------------------------------- NO CLOCK INSERTED -------------------------------------------------------
//    input wire [FP_SIZE-1:0] min_eigen_values [0:MIN_PC_NUM-1],
//    input wire [FP_SIZE-1:0] min_principal_comps [0:MIN_PC_NUM-1],
//    output wire [FP_SIZE-1:0] min_pc_score
//------------------------------------------------------------------------------------------------------------------------
//****************************************************************************************************************************************************
//********************************************************* USING FLOATING POINT *********************************************************************
//---------------------------------------------- CLOCK INSERTED ----------------------------------------------------------
//    input wire clk, reset,
//    input real min_eigen_values [0:MIN_PC_NUM-1],
//    input real min_principal_comps [0:MIN_PC_NUM-1],
//    output real min_pc_score
// -----------------------------------------------------------------------------------------------------------------------
//---------------------------------------------- NO CLOCK INSERTED -------------------------------------------------------
    input real min_eigen_values [0:MIN_PC_NUM-1],
    input real min_principal_comps [0:MIN_PC_NUM-1],
    output real min_pc_score
//------------------------------------------------------------------------------------------------------------------------

//***************************************************************************************************************************************************

);

//********************************************************* USING 64 BIT BINARY *********************************************************************

//-------------------------------------------- NO CLOKC INSERTED -------------------------------------------------------
//wire [FP_SIZE-1:0] temp [0:PC_NUM-1];
//wire [FP_SIZE-1:0] sum_sq;

// assign sum_sq = {FP_SIZE{1'b0}};
//genvar i;
//generate
//    for (i = 0; i < PC_NUM; i = i + 1) begin : SQ_LOOP
//        assign temp[i] = min_principal_comps[i] * min_principal_comps[i] / min_eigen_values[i];
//        assign sum_sq = sum_sq + temp[i];
//    end
//endgenerate
//------------------------------------------------------------------------------------------------------------------------

//---------------------------------------------- CLOCK INSERTED ----------------------------------------------------------
//reg [FP_SIZE-1:0] temp [0:PC_NUM-1];
//reg [FP_SIZE-1:0] sum_sq;

//always @(*) begin
//    if (reset) begin
//        sum_sq <= {FP_SIZE{1'b0}};
//    end else begin
//        sum_sq <= {FP_SIZE{1'b0}};
//        for (int i = 0; i < MIN_PC_NUM; i = i + 1) begin
//            temp[i] <= min_principal_comps[i] * min_principal_comps[i] / min_eigen_values[i];
//            sum_sq <= sum_sq + temp[i];
//        end
//    end
//end
//------------------------------------------------------------------------------------------------------------------------

//****************************************************************************************************************************************************


//********************************************************* USING FLOATING POINT *********************************************************************

//-------------------------------------------- NO CLOKC INSERTED -------------------------------------------------------
    integer i;
    real sum_sq;
//    real POS_INF = $bitstoreal(32'h7f800000); // Positive infinity
//    real NEG_INF = $bitstoreal(32'hff800000); // Negative infinity
    always @(*) begin
        sum_sq = 0;
        for (i = 0; i < MIN_PC_NUM; i = i + 1) begin
            sum_sq = sum_sq + ((min_principal_comps[i] * min_principal_comps[i]) / min_eigen_values[i]);
        end
    end

// assign sum_sq = 0;
//genvar i;
//generate
//    for (i = 0; i < MIN_PC_NUM; i = i + 1) begin : SQ_LOOP
//        assign temp[i] = (min_principal_comps[i] * min_principal_comps[i]) / min_eigen_values[i];
//        assign sum_sq = sum_sq + temp[i];
//    end

//for (i = 0; i < MIN_PC_NUM; i = i + 1) begin : SQ_LOOP
//    if (min_eigen_values[i] != 0) begin
//        temp[i] = (min_principal_comps[i] * min_principal_comps[i]) / min_eigen_values[i];
//        if (!$isinf(temp[i]) && !$isnan(temp[i])) begin
//            sum_sq = sum_sq + temp[i];
//        end
//    end else begin
//        // Handle division by zero
//        temp[i] = 0;
//    end
//end

//endgenerate

//initial begin
//        sum_sq = 0;
//        for (int i = 0; i < MIN_PC_NUM; i = i + 1) begin
//            if (min_eigen_values[i] != 0) begin
//                temp[i] = (min_principal_comps[i] * min_principal_comps[i]) / min_eigen_values[i];
//                if (temp[i] == POS_INF || temp[i] == NEG_INF) begin
//                    temp[i] = 0; // Handle infinity
//                end
//                sum_sq = sum_sq + temp[i];
//            end else begin
//                // Handle division by zero
//                temp[i] = 0;
//            end
//        end
//        min_pc_score = sum_sq;
//    end
//------------------------------------------------------------------------------------------------------------------------

//---------------------------------------------- CLOCK INSERTED ----------------------------------------------------------
//real temp [0:PC_NUM-1];
//real sum_sq;

//always @(*) begin
//    if (reset) begin
//        sum_sq <= 0;
//    end else begin
//        sum_sq <= 0;
//        for (int i = 0; i < MIN_PC_NUM; i = i + 1) begin
//            temp[i] <= min_principal_comps[i] * min_principal_comps[i] / min_eigen_values[i];
//            sum_sq <= sum_sq + temp[i];
//        end
//    end
//end

//------------------------------------------------------------------------------------------------------------------------

//****************************************************************************************************************************************************

assign min_pc_score = sum_sq;

endmodule
