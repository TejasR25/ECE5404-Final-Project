//`timescale 1ns / 1ps
//       file_sample_input = $fopen("train_sample.txt", "r");
//       if (file_sample_input == 0) begin
//       $display("FILE IS NULL");
//       $finish;
      // end
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.05.2024 09:28:12
// Design Name: 
// Module Name: nsl_ids_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module nsl_ids_tb;
//Parameters
    parameter PC_NUM = 32, MAJ_PC_NUM = 10,MIN_PC_NUM = 5, FP_SIZE = 64;
        
        // Inputs and Outputs
   // logic clk;
   // logic reset;
    reg [FP_SIZE-1:0] sorted_eigen_values [0:PC_NUM -1];
    reg [FP_SIZE-1:0] sorted_eigen_vectors [0:PC_NUM-1][0:PC_NUM-1];
    reg [FP_SIZE-1:0] input_samples [0:PC_NUM -1];
    logic ids_out;
    //logic ids_out_f;
    
    //Instatiating the DUT
    nsl_ids #(.PC_NUM(PC_NUM), .MAJ_PC_NUM(MAJ_PC_NUM), .MIN_PC_NUM(MIN_PC_NUM), .FP_SIZE(FP_SIZE))
    dut(
      //  .clk(clk), .reset(reset),
        .sorted_eigen_values(sorted_eigen_values),   // Defining an array made up of (PC_NUM) elements each of (FP_SIZE) bits
        .sorted_eigen_vectors(sorted_eigen_vectors), // Defining an array made up of (PC_NUM * PC_NUM) elements each of (FP_SIZE) bits
        .input_samples(input_samples),               // Defining an array made up of (PC_NUM) elements each of (FP_SIZE) bits 
        .ids_out(ids_out)
    );
    
//    // Read data from CSV file and apply it to inputs
//   initial begin
   
//       // Variables for reading CSV file
//       integer file_eigen_values;
//       integer file_eigen_vectors;
//       integer file_sample_input;
       
//       bit [FP_SIZE-1:0] eigen_value_dec;
//       bit [FP_SIZE-1:0] eigen_vector_dec;
//       bit [FP_SIZE-1:0] sample_input_dec;

//       // Open the CSV files for reading 
//       file_eigen_values = $fopen("\Post PCA inputs\sorted_eig_val", "r");
//       file_eigen_vectors = $fopen("\Post PCA inputs\sorted_eig_vec", "r");
//       file_sample_input = $fopen("\Post PCA inputs\train_sample", "r");
       
//       // Read input samples
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           $fscanf(file_sample_input, "%d,", sample_input_dec);
//           input_samples[i] = $bitstoreal(sample_input_dec);
//       end
       
//       // Read sorted eigen values
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           $fscanf(file_eigen_values, "%d,", eigen_value_dec);
//           sorted_eigen_values[i] = $bitstoreal(eigen_value_dec);
//       end

//       // Read sorted eigen vectors
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           for (int j = 0; j < PC_NUM; j = j + 1) begin
//               $fscanf(file_eigen_vectors, "%d,", eigen_vector_dec);
//               sorted_eigen_vectors[i][j] = $bitstoreal(eigen_vector_dec);
//           end
//       end

//       // Close the CSV files
//       $fclose(file_eigen_values);
//       $fclose(file_eigen_vectors);
//       $fclose(file_sample_input);
       
//timeunit 1ns;

//timeprecision 100ps;
       
       // Read eigen_values  data from file
   initial begin
   
   //ids_out_f = 1'b0;
    // Repeat for all PC_NUM * PC_NUM elements

  $display($time, " << Starting the Simulation >>");
  //  reset = 1'b1;
   // clk = 1;
//begin
//#5 reset = ~reset;
//end

//begin forever
//#5 clk = ~clk; // Toggle the clock every 5 time units 
//end   
//       integer file_sample_input;
//       integer file_eigen_values;
//       integer file_eigen_vectors;
       
//       real sample_input_dec;
//       real sorted_eigen_value_dec;
//       real sorted_eigen_vector_dec;
       
//       file_sample_input = $fopen("train_sample.csv", "r");
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           $fscanf(file_sample_input, "%d,", sample_input_dec);
//           input_samples[i] = $realtobits(sample_input_dec);
//       end
//       $fclose(file_sample_input); 
         

//       file_eigen_values = $fopen("sorted_eig_val.csv", "r");
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           $fscanf(file_eigen_values, "%d\n", sorted_eigen_value_dec);
//           sorted_eigen_values[i] = $realtobits(sorted_eigen_value_dec);
//       end
//       $fclose(file_eigen_values);

//       // Read long_vector data from file
//       file_eigen_vectors = $fopen("sorted_eig_vec.csv", "r");
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           for (int j = 0; j < PC_NUM; j = j + 1) begin
//               $fscanf(file_eigen_vectors, "%d,", sorted_eigen_vector_dec);
//               sorted_eigen_vectors[i][j] = $realtobits(sorted_eigen_vector_dec);
//           end
//           // Skip the newline character at the end of each line
//           $fgetc(file_eigen_vectors);
//       end
//       $fclose(file_eigen_vectors);
      
      // Manually input values for input_samples
//    input_samples[0] = 64'b;
//    input_samples[1] = 64'b;
    // Repeat for all PC_NUM elements
input_samples[0] = 64'b1011111111000000100010101111011111000100001100011010011011011010;
input_samples[1] = 64'b1011111110100000000101010001110001001000110101101010000110100101;
input_samples[2] = 64'b1011111110110000111011101000111011000010011101101111011000001011;
input_samples[3] = 64'b1011111110000001101001011100011011111001001011011001001110110101;
input_samples[4] = 64'b1011111110111001100101001001001111000000001110110111000011110010;
input_samples[5] = 64'b1011111110011100100101001000000110100011010011001100011111110111;
input_samples[6] = 64'b1011111110001111101101110110001100000011101101010101110010110011;
input_samples[7] = 64'b1011111110100111000111011110000101100011110111100001010111111101;
input_samples[8] = 64'b1011111110100001000001101100001000101011101001110101000110110000;
input_samples[9] = 64'b1011111110010001010001100110100011101100110100101111111101000100;
input_samples[10] = 64'b1011111110100001100000011110110111001010010110011000001101110001;
input_samples[11] = 64'b1011111110011000000111111100011110001010010010110001110110010011;
input_samples[12] = 64'b1011111110101100011010110010010001110000001100000111011001011011;
input_samples[13] = 64'b0011111111111101001010100111111010101011000010100010101010000101;
input_samples[14] = 64'b1011111111000010011110010011000001011100000110000101010110000111;
input_samples[15] = 64'b1011111111000010010000101111010001001111110011101010010001100001;
input_samples[16] = 64'b1011111111000001111001010110001100001110011110111101101111001110;
input_samples[17] = 64'b0100000000010010110101100000011011000110001011101100010111110011;
input_samples[18] = 64'b0100000000010010111001001100011010101100000001110111100101011111;
input_samples[19] = 64'b1100000000010110011011001011011000011100000000000000101000110111;
input_samples[20] = 64'b0011111111001011011011110110111110110001100100100100111000001001;
input_samples[21] = 64'b1011111111011101110000000010111100000000111111101000001000100000;
input_samples[22] = 64'b0011111111110000111010001011110001100011000100111110010011011110;
input_samples[23] = 64'b1011111111111101100101111110011000010011001100000100101101010011;
input_samples[24] = 64'b1100000000000010010100000001100101010100100001011110100101010111;
input_samples[25] = 64'b0011111111001101101111100100011000111110011000100001111101011100;
input_samples[26] = 64'b1011111111011110101000000001000100110001001110100010100110101000;
input_samples[27] = 64'b1011111111011000001011011111101110010010011010110111110000011110;
input_samples[28] = 64'b1011111111000011011000010011010001011111001101001100110011000100;
input_samples[29] = 64'b1011111110111011100110101011111011011001111111000101011101011001;
input_samples[30] = 64'b0100000000010011100001101101010101010000011011000101010001001101;
input_samples[31] = 64'b0100000000010011111000011111111011100010111101111100111010001010;


// Manually input values for sorted_eigen_values
sorted_eigen_values[0] = 64'b0100000000010000000001111111111001010110000100000100000110111001;
sorted_eigen_values[1] = 64'b0100000000001011101110101110010000101010011100010110011001111101;
sorted_eigen_values[2] = 64'b0100000000000110110111110101100001110100100000110000010011011011;
sorted_eigen_values[3] = 64'b0100000000000001010100101100100100000100000010000101000101111100;
sorted_eigen_values[4] = 64'b0011111111111111001110110110001010101100010010111010010101110111;
sorted_eigen_values[5] = 64'b0011111111111000010010001111000110100110000011101111011111001010;
sorted_eigen_values[6] = 64'b0011111111110110000101110101000111110000110110000011110111101000;
sorted_eigen_values[7] = 64'b0011111111110101100001010000101111111100100011001011010011110101;
sorted_eigen_values[8] = 64'b0011111111110011111111001011010100000101001100111101101101101011;
sorted_eigen_values[9] = 64'b0011111111110010001001010111100010111110101110000110101000011101;
sorted_eigen_values[10] = 64'b0011111111110001001101111001011001000011001101111001010100111111;
sorted_eigen_values[11] = 64'b0011111111110000101100011100000001011010100000100100111101010011;
sorted_eigen_values[12] = 64'b0011111111101111111011101011010011011110000110000100101100010010;
sorted_eigen_values[13] = 64'b0011111111101111101011000011001010110101011110111011001001110101;
sorted_eigen_values[14] = 64'b0011111111101101001111001001100111001111110001011000001110010010;
sorted_eigen_values[15] = 64'b0011111111101011011110100100011010100001001111011011011001110110;
sorted_eigen_values[16] = 64'b0011111111100111011000000001001011110110001101010110100011101110;
sorted_eigen_values[17] = 64'b0011111111100100011010011100100001101001000010101110000010011101;
sorted_eigen_values[18] = 64'b0011111111100010101111010101110010011011101000100010001101101100;
sorted_eigen_values[19] = 64'b0011111111100001101100010010110000011000110010000000111110110100;
sorted_eigen_values[20] = 64'b0011111111100001010010111011011010000010011101111001010011000101;
sorted_eigen_values[21] = 64'b0011111111011111001110001001001001000001001010011000101101100010;
sorted_eigen_values[22] = 64'b0011111111011001011110101101100000100001000011100101111110111010;
sorted_eigen_values[23] = 64'b0011111111010001000100011001101110100010001010010110101010100001;
sorted_eigen_values[24] = 64'b0011111111001110110011001010111010110010001001010010100111100011;
sorted_eigen_values[25] = 64'b0011111111000111111110010011101100000111010010011011000111111100;
sorted_eigen_values[26] = 64'b0011111110111111000000111010001010010101111000001110000000111101;
sorted_eigen_values[27] = 64'b0011111110111101100010100001100011000111001111110000011111011010;
sorted_eigen_values[28] = 64'b0011111110111011011101101111101111110111111100111011001110000010;
sorted_eigen_values[29] = 64'b0011111110101100001110010011010010011101010010111001101000100100;
sorted_eigen_values[30] = 64'b0011111110010000101000010001001110010001010000011110000000011101;
sorted_eigen_values[31] = 64'b0011111101000001011011001011100011010011110110000010110000111000;

    // Repeat for all PC_NUM elements

// Manually input values for sorted_eigen_vectors
sorted_eigen_vectors[0][0] = 64'b1011111110011011101010111100100011011011011001000101001110000100;
sorted_eigen_vectors[0][1] = 64'b1011111111010001110011001101111110101000001010111100000010011001;
sorted_eigen_vectors[0][2] = 64'b1011111110100110101111111001110111110101100000101000111001011111;
sorted_eigen_vectors[0][3] = 64'b1011111110111100001010011111001000000100001001001110100101100110;
sorted_eigen_vectors[0][4] = 64'b0011111110110101011011111000111100010101110110110100011001100001;
sorted_eigen_vectors[0][5] = 64'b0011111111010010100010010010110001101100011010001010001011000001;
sorted_eigen_vectors[0][6] = 64'b0011111111000000110010111100001111001001010010000000001101100011;
sorted_eigen_vectors[0][7] = 64'b0011111101110011101000010111000011010000011001101001101011110100;
sorted_eigen_vectors[0][8] = 64'b0011111110101000101000110010001101001110100101110001110101110101;
sorted_eigen_vectors[0][9] = 64'b1011111111001010001011111000100100000100010000001100101100101011;
sorted_eigen_vectors[0][10] = 64'b1011111111001011111100010000110010101110100001010110101110001001;
sorted_eigen_vectors[0][11] = 64'b0011111111010100101111101011101011000100101101110110110011010010;
sorted_eigen_vectors[0][12] = 64'b0011111111000010111010001011110000110100101001001111111001111110;
sorted_eigen_vectors[0][13] = 64'b0011111110010110100001001101010011110000110101100110111101111110;
sorted_eigen_vectors[0][14] = 64'b0011111110001110000001000111001010110000010111001010010100101001;
sorted_eigen_vectors[0][15] = 64'b1011111110010101101001110010001101110011101100010100001101110110;
sorted_eigen_vectors[0][16] = 64'b1011111110111100001111010011001110001011101100001111101110100101;
sorted_eigen_vectors[0][17] = 64'b0011111111001110111110001101010101101000011001100011101010011001;
sorted_eigen_vectors[0][18] = 64'b1011111111011000110110111101011001011110010001001110011111100110;
sorted_eigen_vectors[0][19] = 64'b0011111111010001111110011100101011110000001110110001111100011010;
sorted_eigen_vectors[0][20] = 64'b1011111111000011000110010000010111000000000100011101110100100100;
sorted_eigen_vectors[0][21] = 64'b0011111111010110000101001000101000100101000111011011010001110000;
sorted_eigen_vectors[0][22] = 64'b1011111111010101011110010001101011011110001011110001000100010000;
sorted_eigen_vectors[0][23] = 64'b0011111110111001011101110001100111001111100101010100110011000100;
sorted_eigen_vectors[0][24] = 64'b1011111110001011100010010101110001010110010000110101101101100001;
sorted_eigen_vectors[0][25] = 64'b1011111110110111110101001011110101000111001000101000111000011111;
sorted_eigen_vectors[0][26] = 64'b1011111110101101101010000001001000110001000010110011011010010010;
sorted_eigen_vectors[0][27] = 64'b1011111110001001010101101101110110100011101110100001110011110001;
sorted_eigen_vectors[0][28] = 64'b1011111110101101001000111001000111000010011001110010110010000010;
sorted_eigen_vectors[0][29] = 64'b0011111100010011110010101000111110011001001001111101011111100100;
sorted_eigen_vectors[0][30] = 64'b0011111101110100001010011000000011111001101110011011001111110101;
sorted_eigen_vectors[0][31] = 64'b0011111101001001110000111010100011110001011001110011010100110000;
sorted_eigen_vectors[1][0] = 64'b0011111101100101100001010010110001010010001001110010110111001001;
sorted_eigen_vectors[1][1] = 64'b1011111110100001001111011001001000110001111001010101011111111111;
sorted_eigen_vectors[1][2] = 64'b1011111101111100110100110011101010110010110010100100111011111001;
sorted_eigen_vectors[1][3] = 64'b0011111110010011110110100100111010100000011000110101000110001000;
sorted_eigen_vectors[1][4] = 64'b1011111100111101101000010001000001110011011100110001011101111000;
sorted_eigen_vectors[1][5] = 64'b0011111111000001110100101111001101110001111011101001010100100101;
sorted_eigen_vectors[1][6] = 64'b1011111111100011111101010100010010111100000100101110000010010001;
sorted_eigen_vectors[1][7] = 64'b0011111111001111010110000001000010010010110000100101111010111000;
sorted_eigen_vectors[1][8] = 64'b0011111111000010001001101010011101111000001100011100000100110011;
sorted_eigen_vectors[1][9] = 64'b1011111111000100111111101011011111001001101110110111011000010100;
sorted_eigen_vectors[1][10] = 64'b0011111110101000001110010010001110010100110100011111111110011001;
sorted_eigen_vectors[1][11] = 64'b0011111110101001010110101000001111010001100100010111110100101111;
sorted_eigen_vectors[1][12] = 64'b0011111110010111110000100111011101101001110001110100011100101110;
sorted_eigen_vectors[1][13] = 64'b1011111110001011010001110010110100101101000111111100100110101110;
sorted_eigen_vectors[1][14] = 64'b1011111110110011101110111000101001000001001100011110001000010100;
sorted_eigen_vectors[1][15] = 64'b0011111110101101110100011011101001011011101010101000010101101001;
sorted_eigen_vectors[1][16] = 64'b0011111111000100100001111100000010111101010011011100101101111011;
sorted_eigen_vectors[1][17] = 64'b1011111111011011001011000010001111111001110000000001000110011110;
sorted_eigen_vectors[1][18] = 64'b1011111110010001100000110111000111000111110010111100001001010100;
sorted_eigen_vectors[1][19] = 64'b0011111111100000000011001101111111000011111110001001010111101000;
sorted_eigen_vectors[1][20] = 64'b0011111110110100011001010001101010110110010001010001111100001010;
sorted_eigen_vectors[1][21] = 64'b1011111110101000010011001001111110011001001001101010110001011100;
sorted_eigen_vectors[1][22] = 64'b0011111110100101000010110000000101010101110001010000110110110011;
sorted_eigen_vectors[1][23] = 64'b0011111110000001001110010010010110010110001110001001111110101110;
sorted_eigen_vectors[1][24] = 64'b0011111110000101010110010010110010000000100100000110010100000110;
sorted_eigen_vectors[1][25] = 64'b1011111101010110111011011111001101110000011111101111001101001001;
sorted_eigen_vectors[1][26] = 64'b0011111101000111011101100001010010001111101100011011001100111001;
sorted_eigen_vectors[1][27] = 64'b0011111101011000101010101110101000100110010010001010010010001011;
sorted_eigen_vectors[1][28] = 64'b1011111101101110101010111001101110111011010110100101100011010111;
sorted_eigen_vectors[1][29] = 64'b1011111100110001110000101100101110100110010110100011111111000110;
sorted_eigen_vectors[1][30] = 64'b1011111100100110100101000101111000111101010010000001011001110110;
sorted_eigen_vectors[1][31] = 64'b0011111100110110100001001111111010101111001001101011101101010100;
sorted_eigen_vectors[2][0] = 64'b0011111101100000111100001000011110110100111001111101000011110010;
sorted_eigen_vectors[2][1] = 64'b1011111110110001100010011101001011101010111101111000110001111110;
sorted_eigen_vectors[2][2] = 64'b1011111110111010110001110011010010111100011111110101000111000010;
sorted_eigen_vectors[2][3] = 64'b0011111110101100011110000101100010000110111000011001111001101001;
sorted_eigen_vectors[2][4] = 64'b0011111110001110010000001001100101111010101111000000001100100000;
sorted_eigen_vectors[2][5] = 64'b0011111111000010100000100000111001111010110110010011100101100101;
sorted_eigen_vectors[2][6] = 64'b1011111111100100000110011101010100100100100000101001001100110111;
sorted_eigen_vectors[2][7] = 64'b0011111111000111101000100010011100110100000010011110101000011001;
sorted_eigen_vectors[2][8] = 64'b0011111110111011100011010011000010110101101011000011111111000110;
sorted_eigen_vectors[2][9] = 64'b1011111110110010010110101110011110011001101010110011010001111000;
sorted_eigen_vectors[2][10] = 64'b1011111110010000011101001100010000011110011111100001011100111001;
sorted_eigen_vectors[2][11] = 64'b0011111101111000111101011010010100100010110111001100000101010001;
sorted_eigen_vectors[2][12] = 64'b0011111110001001110011010001111111001001011101001101110100100101;
sorted_eigen_vectors[2][13] = 64'b0011111110001001100100001000010000111111010110000110001100110101;
sorted_eigen_vectors[2][14] = 64'b1011111110000000101101111010000100001000111100110100110110100111;
sorted_eigen_vectors[2][15] = 64'b1011111110011110001111100111110010110000100001100100000110110100;
sorted_eigen_vectors[2][16] = 64'b1011111111000100011001111010100110101000101010010000101000110110;
sorted_eigen_vectors[2][17] = 64'b0011111111011001011011011111010111001000110101100011000100011111;
sorted_eigen_vectors[2][18] = 64'b1011111110001011101100010110011100111110101011010101011001010010;
sorted_eigen_vectors[2][19] = 64'b1011111111100001111010100010110110001111100001110111001010100111;
sorted_eigen_vectors[2][20] = 64'b1011111110111110111100000100111000001110101001011010010101100010;
sorted_eigen_vectors[2][21] = 64'b0011111110011010111111000011011011010011110100010001111000100110;
sorted_eigen_vectors[2][22] = 64'b1011111110010101111001101001000000000101110101001011011000011010;
sorted_eigen_vectors[2][23] = 64'b1011111110010100000010111111001101111011100011001000111010010101;
sorted_eigen_vectors[2][24] = 64'b1011111101111001101111100000110001111001101111010100111111110001;
sorted_eigen_vectors[2][25] = 64'b0011111110000100000000110111110000110000001010011101101111111000;
sorted_eigen_vectors[2][26] = 64'b0011111101110101110101000111000010111110111111111010001011000111;
sorted_eigen_vectors[2][27] = 64'b1011111101100110101101011011011010001100101111111110010011010111;
sorted_eigen_vectors[2][28] = 64'b0011111101010010100000000000101011001000010111110011011110000100;
sorted_eigen_vectors[2][29] = 64'b1011111101001000010110000001011010111101100100010000000110010011;
sorted_eigen_vectors[2][30] = 64'b0011111100110011110101000011111101110011001100100011101010011010;
sorted_eigen_vectors[2][31] = 64'b1011111101010001101111110011001001101110011011011110101100001000;
sorted_eigen_vectors[3][0] = 64'b1011111101100001110000011000101111000111010011101110110101111000;
sorted_eigen_vectors[3][1] = 64'b1011111110100000100100000111000000110111100000111101100110100110;
sorted_eigen_vectors[3][2] = 64'b1011111110101100100101001110100100111110010000110000001100000011;
sorted_eigen_vectors[3][3] = 64'b1011111110000001100100110111111100111010100011110110010010101001;
sorted_eigen_vectors[3][4] = 64'b1011111110000011011110110101000110110010011001011110101100001101;
sorted_eigen_vectors[3][5] = 64'b0011111110101000010111110101010100111110011111000100110010110111;
sorted_eigen_vectors[3][6] = 64'b1011111110100110010001111010111010101010110110011011000001101110;
sorted_eigen_vectors[3][7] = 64'b1011111110110000100001000010110110000000010110001111001101111000;
sorted_eigen_vectors[3][8] = 64'b0011111111001100011000001101100110011110010111010111111101001011;
sorted_eigen_vectors[3][9] = 64'b0011111111100011011010100010110101010110100000111000111111001101;
sorted_eigen_vectors[3][10] = 64'b1011111111001011100110100010111111000010101111010100010110010100;
sorted_eigen_vectors[3][11] = 64'b0011111110111010011111100010100110101001101111011100101100111000;
sorted_eigen_vectors[3][12] = 64'b0011111110100100011101100011000110110110110000101111000010011110;
sorted_eigen_vectors[3][13] = 64'b1011111110010010110100100010010010001101000101100101011000001010;
sorted_eigen_vectors[3][14] = 64'b1011111111000011101111011011100100011101110111111101001111101101;
sorted_eigen_vectors[3][15] = 64'b0011111111100101110110001111110110001000111000101101010100010000;
sorted_eigen_vectors[3][16] = 64'b1011111110010100010111010010101001110100010111100111000010000111;
sorted_eigen_vectors[3][17] = 64'b1011111110101101000010111001100010011111001110110010000110000011;
sorted_eigen_vectors[3][18] = 64'b1011111110111011000111011101100011010000011001000011001010101011;
sorted_eigen_vectors[3][19] = 64'b1011111110100111101011010100001100101011110101111100001111100101;
sorted_eigen_vectors[3][20] = 64'b0011111110011000011101100001011011100101100000101010101111100001;
sorted_eigen_vectors[3][21] = 64'b0011111110011000001000010011010101000001101010110010001111101000;
sorted_eigen_vectors[3][22] = 64'b0011111101111111000101010010101011011011110000100111101100010001;
sorted_eigen_vectors[3][23] = 64'b0011111110101011010010000110110110100110101011110111111111010010;
sorted_eigen_vectors[3][24] = 64'b1011111101011111001110101000100110100100101110011011110100000011;
sorted_eigen_vectors[3][25] = 64'b1011111101110011110001000000101111011001000110111010010001100000;
sorted_eigen_vectors[3][26] = 64'b1011111101011100110000110100000111001001010000111111000110001100;
sorted_eigen_vectors[3][27] = 64'b1011111100110011011000000111110010011000101100000010101010101001;
sorted_eigen_vectors[3][28] = 64'b1011111101001111100100010101110001001000111101110000011000101101;
sorted_eigen_vectors[3][29] = 64'b1011111100110011110101010111100100011000010100100101001000110010;
sorted_eigen_vectors[3][30] = 64'b0011111101000001011110110101111001011100110010111001111010110000;
sorted_eigen_vectors[3][31] = 64'b1011111101100000101101000001101001010000001110101001101011010001;
sorted_eigen_vectors[4][0] = 64'b0011111110000010010101100110111010010000101101100110001101100000;
sorted_eigen_vectors[4][1] = 64'b1011111110110000110001111000011111010110110000001000010011110001;
sorted_eigen_vectors[4][2] = 64'b0011111110100100001010100111100101101111000001100001101000101100;
sorted_eigen_vectors[4][3] = 64'b0011111100110011111011011011111010111011011110110100110101011010;
sorted_eigen_vectors[4][4] = 64'b1011111110011100010010001100101110011001001010000100010110011000;
sorted_eigen_vectors[4][5] = 64'b0011111110110000100110101101011111101100011110100011111010100111;
sorted_eigen_vectors[4][6] = 64'b1011111110001110000110111010110000101011011101110001010100001100;
sorted_eigen_vectors[4][7] = 64'b1011111110011010010001110101011101011101011111100010011110110000;
sorted_eigen_vectors[4][8] = 64'b1011111111000011011101001011110010011011101101011001001000001111;
sorted_eigen_vectors[4][9] = 64'b0011111111001101110011010010101110111110011101100000110011000100;
sorted_eigen_vectors[4][10] = 64'b0011111111100110010011110110100110000101111110011000100011110001;
sorted_eigen_vectors[4][11] = 64'b0011111111000110100101101010111111110000111010101111011101101101;
sorted_eigen_vectors[4][12] = 64'b0011111111001010110011010100111100100011100000101101111011111011;
sorted_eigen_vectors[4][13] = 64'b0011111111010101101110100001001000100110101011000111100100000001;
sorted_eigen_vectors[4][14] = 64'b1011111111001011010110010011010000110101010110111100101110000001;
sorted_eigen_vectors[4][15] = 64'b1011111110101000011111101101000001011110101010000001000110010111;
sorted_eigen_vectors[4][16] = 64'b1011111111010110001101100001011101010000000010000111100101110000;
sorted_eigen_vectors[4][17] = 64'b1011111110010010000100001110100100111000000001000001010011111000;
sorted_eigen_vectors[4][18] = 64'b1011111111000101101111001110011001101110101110011100101101100000;
sorted_eigen_vectors[4][19] = 64'b0011111110110011000010101110101111000010000001101010101101000111;
sorted_eigen_vectors[4][20] = 64'b1011111110111110001011101110001010100011011111100000000000110101;
sorted_eigen_vectors[4][21] = 64'b1011111111000000000100000001111011110011101000011100010110101110;
sorted_eigen_vectors[4][22] = 64'b0011111110100000001101101001010000011110111110110001110010011100;
sorted_eigen_vectors[4][23] = 64'b1011111101110100100001010101110000000100000101011110000100100010;
sorted_eigen_vectors[4][24] = 64'b0011111110011010110101100011001011011100010001110101010100000101;
sorted_eigen_vectors[4][25] = 64'b0011111110000011001101000100100011110000010011110010110011011001;
sorted_eigen_vectors[4][26] = 64'b1011111101010011111100000001101111000011011111110110111111111010;
sorted_eigen_vectors[4][27] = 64'b1011111110000001110111011100011011110000011111100001100110101001;
sorted_eigen_vectors[4][28] = 64'b1011111101000101111100100111011110010110010100100011110000100011;
sorted_eigen_vectors[4][29] = 64'b1011111101010100101010010010001010010011110110100101110100100010;
sorted_eigen_vectors[4][30] = 64'b1011111101000101010111000010100100100100110110100100101001000000;
sorted_eigen_vectors[4][31] = 64'b1011111100110111000100100010100110101000001101000110001000101111;
sorted_eigen_vectors[5][0] = 64'b1011111101110110101000100100100001100010101010000111011000000000;
sorted_eigen_vectors[5][1] = 64'b1011111110101000000010000011100101010111101011100110110111001101;
sorted_eigen_vectors[5][2] = 64'b1011111110100010000110001111110010111101100011110010001011011100;
sorted_eigen_vectors[5][3] = 64'b0011111101101111010110011001110100110011101100001000010111101111;
sorted_eigen_vectors[5][4] = 64'b0011111110000101111000011110111010100001110000101001001011101111;
sorted_eigen_vectors[5][5] = 64'b0011111110110110010010000111010110101101111001001011111100111001;
sorted_eigen_vectors[5][6] = 64'b1011111110111010100111101110100110110111000001111010111110111110;
sorted_eigen_vectors[5][7] = 64'b1011111110110011001001000110110100010100010101011101111111001100;
sorted_eigen_vectors[5][8] = 64'b0011111111000100001001000000111000001010100100010001001101111000;
sorted_eigen_vectors[5][9] = 64'b0011111111100011010111010100111110000001111111100101111011001110;
sorted_eigen_vectors[5][10] = 64'b1011111111001100001111110101000011110100001110111101000011110100;
sorted_eigen_vectors[5][11] = 64'b0011111111000001000100000011010111100101010010001000110111100011;
sorted_eigen_vectors[5][12] = 64'b0011111101011010110001011110001100000101101010111011100001000101;
sorted_eigen_vectors[5][13] = 64'b1011111110101110101110001110000111100111010101110101101001010111;
sorted_eigen_vectors[5][14] = 64'b0011111111000010011010101011101110001100110000001000001010001110;
sorted_eigen_vectors[5][15] = 64'b1011111111100101111011110010110110011101001101001011010000101010;
sorted_eigen_vectors[5][16] = 64'b0011111101011110010100000110000001001111000010100100100101001110;
sorted_eigen_vectors[5][17] = 64'b1011111110111001101101111001000011101110111111001110110101110110;
sorted_eigen_vectors[5][18] = 64'b1011111110100100001010100001001100101101010011011010100100111000;
sorted_eigen_vectors[5][19] = 64'b0011111110100111110110101100000111010011011011001100000000100101;
sorted_eigen_vectors[5][20] = 64'b1011111110000101101101001101101000101110000100010101010111010111;
sorted_eigen_vectors[5][21] = 64'b1011111110110000001001001101110110000001110010100000000100110000;
sorted_eigen_vectors[5][22] = 64'b0011111110010011111001110010101100011000010011000110110111111001;
sorted_eigen_vectors[5][23] = 64'b0011111110101000111100010100011101000100001011011100001001111111;
sorted_eigen_vectors[5][24] = 64'b0011111101110101010011010011000111111001010000010010000111010000;
sorted_eigen_vectors[5][25] = 64'b1011111110000101111100111111001011110000100000011001010110000110;
sorted_eigen_vectors[5][26] = 64'b0011111101100010110010000010011101101100001110111010000011101110;
sorted_eigen_vectors[5][27] = 64'b1011111101110110111101001111000111111010110000001011010111110101;
sorted_eigen_vectors[5][28] = 64'b0011111100110110110011000100111010011100111011101000111100100110;
sorted_eigen_vectors[5][29] = 64'b0011111100101110010011101010111100110111000000111001100101010101;
sorted_eigen_vectors[5][30] = 64'b1011111100111001111101001010001110001001110000000001010001100000;
sorted_eigen_vectors[5][31] = 64'b1011111101011101000110010001001001111011111000100000100111000011;
sorted_eigen_vectors[6][0] = 64'b1011111110000000101100000111110001010010000010010001000111001011;
sorted_eigen_vectors[6][1] = 64'b1011111111000110010101010001100001000111001001110110001001110011;
sorted_eigen_vectors[6][2] = 64'b1011111111011010010000011100111011001011110110010000001111101011;
sorted_eigen_vectors[6][3] = 64'b1011111110111000100101000111101101111000111111100010110111011001;
sorted_eigen_vectors[6][4] = 64'b1011111110110110111100000001110001010000001011000101100101110111;
sorted_eigen_vectors[6][5] = 64'b1011111111001110101100010110111110110011011011100011011011111001;
sorted_eigen_vectors[6][6] = 64'b1011111110010100001110010011000111101111010101101100010000110110;
sorted_eigen_vectors[6][7] = 64'b0011111111010000000001110011100010111110010001000110110101100000;
sorted_eigen_vectors[6][8] = 64'b1011111111011000000101001111100010111011000100111101010110110100;
sorted_eigen_vectors[6][9] = 64'b0011111110110110101010011101101110110000110001100110011100100101;
sorted_eigen_vectors[6][10] = 64'b1011111110111011101000110100010000000011010011001011110010101011;
sorted_eigen_vectors[6][11] = 64'b0011111110011000101111100101011100011000110110000100111110001100;
sorted_eigen_vectors[6][12] = 64'b0011111110101000111100011010010110011110101010111010101011101111;
sorted_eigen_vectors[6][13] = 64'b0011111110010100110110001011101011100000000100111001101111100011;
sorted_eigen_vectors[6][14] = 64'b1011111110000011110111111011000001001000100100001000010000010000;
sorted_eigen_vectors[6][15] = 64'b0011111101111000101111000110101011110010001001011100110111010010;
sorted_eigen_vectors[6][16] = 64'b1011111101000000011110100110111100010111011011010111011111010001;
sorted_eigen_vectors[6][17] = 64'b0011111110001001111000000011110001010110101111010111110001010010;
sorted_eigen_vectors[6][18] = 64'b0011111110100100000001111100111010001001001101011100010001010010;
sorted_eigen_vectors[6][19] = 64'b0011111110101011010000101100111110100001111010101000001000100110;
sorted_eigen_vectors[6][20] = 64'b0011111101110100000010111111101101100111101001101011100100110101;
sorted_eigen_vectors[6][21] = 64'b1011111110001101001011100111110101001101110010000101111010001101;
sorted_eigen_vectors[6][22] = 64'b0011111110000101101000110011010000101111011111011100001000111001;
sorted_eigen_vectors[6][23] = 64'b0011111110100100000001010110000010110101010100111010101111010001;
sorted_eigen_vectors[6][24] = 64'b1011111100111100010111001010100111111010111010010011100001110111;
sorted_eigen_vectors[6][25] = 64'b1011111101011110111000110010111100110001000100111110011100110101;
sorted_eigen_vectors[6][26] = 64'b0011111100110010000110111001000000110101001111111010011100000011;
sorted_eigen_vectors[6][27] = 64'b1011111100010101101101101110100000001110100001100101000011011011;
sorted_eigen_vectors[6][28] = 64'b0011111101000011010110100010000010011001000101011010010100000010;
sorted_eigen_vectors[6][29] = 64'b0011111100111010010101010000011011001001001111000001101000110000;
sorted_eigen_vectors[6][30] = 64'b1011111101010111011011011101010000011111101011001110101010011001;
sorted_eigen_vectors[6][31] = 64'b0011111111100110011101000000110101010111111110100111110011101111;
sorted_eigen_vectors[7][0] = 64'b1011111110000111000110100001010101011001001010000000001000100010;
sorted_eigen_vectors[7][1] = 64'b1011111111000110000011001001010000111011011010110111010001001011;
sorted_eigen_vectors[7][2] = 64'b1011111111010101111110111110100000011001000101111000110101000001;
sorted_eigen_vectors[7][3] = 64'b1011111110011001010101000110001110001000101000111000110100110001;
sorted_eigen_vectors[7][4] = 64'b1011111110010000110011001010010111100011100001010100111111000010;
sorted_eigen_vectors[7][5] = 64'b0011111110101110111100001101011101111101001001100111010101100000;
sorted_eigen_vectors[7][6] = 64'b0011111110100100100110111101010000101110011001101100100111010101;
sorted_eigen_vectors[7][7] = 64'b1011111111001001100110100011101101011001110111000001101000101000;
sorted_eigen_vectors[7][8] = 64'b0011111111010111000010110011011111010111011110110000001000001000;
sorted_eigen_vectors[7][9] = 64'b1011111110101010100010111110010100000110010110100000001011100111;
sorted_eigen_vectors[7][10] = 64'b0011111111000111010001111000011111011010010011001110000000111000;
sorted_eigen_vectors[7][11] = 64'b1011111110111010111010000001111100101101011110100001001000010111;
sorted_eigen_vectors[7][12] = 64'b1011111110101011010110110100011111100100111100101001010100100000;
sorted_eigen_vectors[7][13] = 64'b1011111110100100000111001100000100010001001100100101100100011101;
sorted_eigen_vectors[7][14] = 64'b0011111110011101111000110110010100000010000111000000110110101000;
sorted_eigen_vectors[7][15] = 64'b0011111110010111000000010000100101101000101001100101001100100001;
sorted_eigen_vectors[7][16] = 64'b1011111110110101001000000110010010100111010001111010010100110101;
sorted_eigen_vectors[7][17] = 64'b0011111111001110010001010001101011100000000101111100011010100101;
sorted_eigen_vectors[7][18] = 64'b0011111111011101100010110001110011011111000110111011001010101111;
sorted_eigen_vectors[7][19] = 64'b0011111111001101010101000001110011111111101001000100111011011011;
sorted_eigen_vectors[7][20] = 64'b1011111110111001111111010001101100000111110000000001110111000010;
sorted_eigen_vectors[7][21] = 64'b1011111110110011001011100010111110111000110000111000110011000110;
sorted_eigen_vectors[7][22] = 64'b0011111110110110000011101001101100010010100101100110011111010010;
sorted_eigen_vectors[7][23] = 64'b0011111111100000101000010000110000001111010111111001011011010110;
sorted_eigen_vectors[7][24] = 64'b1011111110010000110110010111000111101110110000101011101100011000;
sorted_eigen_vectors[7][25] = 64'b1011111110100101101111110101000111111111101010110111011010000100;
sorted_eigen_vectors[7][26] = 64'b1011111101110111111000111011100011110001100010000101111110011100;
sorted_eigen_vectors[7][27] = 64'b1011111101100110001011110101100011000011011110000000000000111001;
sorted_eigen_vectors[7][28] = 64'b0011111100110100101100000101110110010010111001101100010110010011;
sorted_eigen_vectors[7][29] = 64'b1011111101100010000101001011000011000101010001001000111110011001;
sorted_eigen_vectors[7][30] = 64'b1011111100110010111101111011100101000110100111010011100111011011;
sorted_eigen_vectors[7][31] = 64'b0011111101011001010011000000001100111111101010100111101111100001;
sorted_eigen_vectors[8][0] = 64'b1011111110001001111010111101100010011101010001011010011111010001;
sorted_eigen_vectors[8][1] = 64'b1011111111001011010000000101001110010111101011000011100110111010;
sorted_eigen_vectors[8][2] = 64'b1011111111011001111010011111110001001000001111111110001101110111;
sorted_eigen_vectors[8][3] = 64'b1011111110100000111100000111000000101101010111101011111011100010;
sorted_eigen_vectors[8][4] = 64'b1011111110000011101001010111001110010010100001101011011010001011;
sorted_eigen_vectors[8][5] = 64'b0011111110100100010101110111010001100110100000101001100011000101;
sorted_eigen_vectors[8][6] = 64'b0011111110101101110110111110000001001011101000110101010100010100;
sorted_eigen_vectors[8][7] = 64'b1011111111000111011100101100001111001111001101000011001001110011;
sorted_eigen_vectors[8][8] = 64'b0011111111010011011000100000000000100111111011100011111010111011;
sorted_eigen_vectors[8][9] = 64'b1011111110010111000001100001001101010110101000101110011110111111;
sorted_eigen_vectors[8][10] = 64'b0011111111000000110110111001111110101000110011000111000001011100;
sorted_eigen_vectors[8][11] = 64'b1011111110101101101000101001010000110111010101011000010001101111;
sorted_eigen_vectors[8][12] = 64'b1011111110110110111110111011010001100000110100111110101000110011;
sorted_eigen_vectors[8][13] = 64'b1011111110100110010111011011010000111011101100001110110000101111;
sorted_eigen_vectors[8][14] = 64'b0011111110100010110010110001101001010000101110100011100011001001;
sorted_eigen_vectors[8][15] = 64'b1011111100101111111011111101100001011110100111001000011000000001;
sorted_eigen_vectors[8][16] = 64'b1011111110011011111101010000001010110001111001110000000100111011;
sorted_eigen_vectors[8][17] = 64'b0011111110010000000111010110010110110011100011011000011011000101;
sorted_eigen_vectors[8][18] = 64'b0011111110101011010101001010110101110011010011000010110100000000;
sorted_eigen_vectors[8][19] = 64'b0011111110110100110001011000010100000110111100011101010001100110;
sorted_eigen_vectors[8][20] = 64'b0011111110001110001100000101001101101001000111110001011101111110;
sorted_eigen_vectors[8][21] = 64'b0011111110000100001110010111011101101100101000001111010110100011;
sorted_eigen_vectors[8][22] = 64'b1011111110101110000100000110101111101010010111111011101000011111;
sorted_eigen_vectors[8][23] = 64'b1011111111101000111001011001111101110101000001100101001000010101;
sorted_eigen_vectors[8][24] = 64'b0011111110011111000101011000111100111011100110010011001011101010;
sorted_eigen_vectors[8][25] = 64'b0011111110110010011010000011011100000110010000101010011000011010;
sorted_eigen_vectors[8][26] = 64'b0011111110010110110101111101110100011001011111000100111100100001;
sorted_eigen_vectors[8][27] = 64'b0011111110001001000011101101010010011000010011000000111000001111;
sorted_eigen_vectors[8][28] = 64'b0011111110000001011100101000011001011101001000101111101101001001;
sorted_eigen_vectors[8][29] = 64'b0011111101101011001111010011101001110100111100111110111001000111;
sorted_eigen_vectors[8][30] = 64'b1011111101101110110000101110001100111110010001000011010000000110;
sorted_eigen_vectors[8][31] = 64'b0011111110001111111111111111101001100010100100001101110100010101;
sorted_eigen_vectors[9][0] = 64'b1011111110000001001111001011101010110111110111010000000101001111;
sorted_eigen_vectors[9][1] = 64'b1011111111000111000010100111001101110101100101100100001011011001;
sorted_eigen_vectors[9][2] = 64'b1011111111011010110111001001100001011100111000001100001011100111;
sorted_eigen_vectors[9][3] = 64'b1011111110111000111110011011001010010111010110010100111111011110;
sorted_eigen_vectors[9][4] = 64'b1011111110110111000110000100001101111011100100101011101101010001;
sorted_eigen_vectors[9][5] = 64'b1011111111001110001010010100001011000100100100111011001111101101;
sorted_eigen_vectors[9][6] = 64'b1011111110001110011100011101100010111010101000111111001011101101;
sorted_eigen_vectors[9][7] = 64'b0011111111001110110001010000110011000001001100011011101101010111;
sorted_eigen_vectors[9][8] = 64'b1011111111010111000010101000111111000111101010011000110010001010;
sorted_eigen_vectors[9][9] = 64'b0011111110110100011011010111010110111110010100001100011001001100;
sorted_eigen_vectors[9][10] = 64'b1011111110111001010010100101010000010000100101111001010110101011;
sorted_eigen_vectors[9][11] = 64'b0011111110010110000001001110010001111100010101101111110001110010;
sorted_eigen_vectors[9][12] = 64'b0011111110100110100111111111100110001010100101000000110101010111;
sorted_eigen_vectors[9][13] = 64'b0011111110010010101111001000101001010010110010011001000110111100;
sorted_eigen_vectors[9][14] = 64'b1011111110000001010001110001010100100001101110101110100011100001;
sorted_eigen_vectors[9][15] = 64'b0011111101110011011100111110011101011010001111000100010011010010;
sorted_eigen_vectors[9][16] = 64'b0011111101100100000111010110011011111011011001111101110011010010;
sorted_eigen_vectors[9][17] = 64'b0011111101101110001110101110001101101001010011101010010100000100;
sorted_eigen_vectors[9][18] = 64'b0011111110100000011111000110000011101110101111000001011000111011;
sorted_eigen_vectors[9][19] = 64'b0011111110101000010010011100000110010000011111000000100101010010;
sorted_eigen_vectors[9][20] = 64'b0011111101111100010000010101101100011111100101100100100010010101;
sorted_eigen_vectors[9][21] = 64'b1011111110001010101011111010011101110010101110101111111111011010;
sorted_eigen_vectors[9][22] = 64'b0011111110000010000100110110010000110100110000110000100111100011;
sorted_eigen_vectors[9][23] = 64'b0011111110011100101000011101001111100100111111101101110101101000;
sorted_eigen_vectors[9][24] = 64'b1011111101001100010110001000101010101111010111100000001111000011;
sorted_eigen_vectors[9][25] = 64'b1011111101011010101100011011111000010101011101101110101000010000;
sorted_eigen_vectors[9][26] = 64'b1011111101011100010100010001011110111010011000010111001100011000;
sorted_eigen_vectors[9][27] = 64'b1011111100111000111010000111111010001000000001001101110011001110;
sorted_eigen_vectors[9][28] = 64'b0011111101100000111001100101100010100000110011001100001011000001;
sorted_eigen_vectors[9][29] = 64'b0011111011010001100101100110000001111001011000111100110110100101;
sorted_eigen_vectors[9][30] = 64'b0011111101001111110010011101011110111101001100111111000000000111;
sorted_eigen_vectors[9][31] = 64'b1011111111100110110010100010110000000111001001100100111100010101;
sorted_eigen_vectors[10][0] = 64'b1011111101110001100110010010001011111101110111001100001111001111;
sorted_eigen_vectors[10][1] = 64'b1011111110110111110011111010101111100101000110110110011101111011;
sorted_eigen_vectors[10][2] = 64'b1011111110100110111010001100100101011110101011100010110101100011;
sorted_eigen_vectors[10][3] = 64'b0011111110101010000100010110001110110111101010110000010011110001;
sorted_eigen_vectors[10][4] = 64'b0011111110111010000110000101000101111100001010110101100011100011;
sorted_eigen_vectors[10][5] = 64'b0011111111010010101101000011010101111011010100110010101100001101;
sorted_eigen_vectors[10][6] = 64'b0011111110100110100001001111010000111001111000111001100011011000;
sorted_eigen_vectors[10][7] = 64'b1011111111001101101110011110111000011010110110000001110110111101;
sorted_eigen_vectors[10][8] = 64'b1011111111000000100110010111000101000101000110011001100110010110;
sorted_eigen_vectors[10][9] = 64'b1011111111000000111011010101000110110100100001101110101011000011;
sorted_eigen_vectors[10][10] = 64'b1011111111010100000000110001010011010001100101010000011010100110;
sorted_eigen_vectors[10][11] = 64'b0011111111000110111010111111100101101000110111011101110110011011;
sorted_eigen_vectors[10][12] = 64'b0011111111011000001111111110101010010100110100010100110001001001;
sorted_eigen_vectors[10][13] = 64'b0011111111010101110000011001000010001001111001100010011101110111;
sorted_eigen_vectors[10][14] = 64'b1011111111011010011110101101011111110100111010100101011010011100;
sorted_eigen_vectors[10][15] = 64'b1011111110110000011101100000111100000100010000100100101110011111;
sorted_eigen_vectors[10][16] = 64'b0011111111001001110110111000011011100000000001011001100111000000;
sorted_eigen_vectors[10][17] = 64'b1011111110110111001111101111110011011111100000011100100001110100;
sorted_eigen_vectors[10][18] = 64'b0011111111010110010101100101100000001010011000000100111011011010;
sorted_eigen_vectors[10][19] = 64'b1011111111000001010100011110001010101101100000111011010011001011;
sorted_eigen_vectors[10][20] = 64'b0011111110000100101010011000011110000100011010100000001101101101;
sorted_eigen_vectors[10][21] = 64'b1011111111000100100100010110011001000111111100101000000010111010;
sorted_eigen_vectors[10][22] = 64'b0011111110111100111010011111001111101010000101011101011101011010;
sorted_eigen_vectors[10][23] = 64'b1011111110110101000010010100010110111001100111100001101101000101;
sorted_eigen_vectors[10][24] = 64'b0011111101100110010010111010110111000111100010000000110011001001;
sorted_eigen_vectors[10][25] = 64'b0011111110100011011000100000000101000101101111000000001100001011;
sorted_eigen_vectors[10][26] = 64'b0011111110010000100110010010011111011010100011101101111011100110;
sorted_eigen_vectors[10][27] = 64'b0011111101100101011000001010000001101001111101011100001000111000;
sorted_eigen_vectors[10][28] = 64'b0011111110001000110101111001111101101101100100101011010011100001;
sorted_eigen_vectors[10][29] = 64'b0011111101001000010110101100111101111010111111011110000010110000;
sorted_eigen_vectors[10][30] = 64'b1011111101011100101010001010101000110111100000100000011101110111;
sorted_eigen_vectors[10][31] = 64'b1011111101011010011101000000000010011100001111111101000000001011;
sorted_eigen_vectors[11][0] = 64'b0011111101011100111010100110010110000110111100000101001010101010;
sorted_eigen_vectors[11][1] = 64'b1011111110010100010101010110101101001100001100001110011000111001;
sorted_eigen_vectors[11][2] = 64'b0011111101111100101011100011001100100000010001110010001011100011;
sorted_eigen_vectors[11][3] = 64'b0011111101011000111100010000001100011001001100001100011110100001;
sorted_eigen_vectors[11][4] = 64'b0011111101110000100000110100110011010001100001010100100000110110;
sorted_eigen_vectors[11][5] = 64'b0011111110011001100011111000111101101011011100011000001000101001;
sorted_eigen_vectors[11][6] = 64'b0011111101100100010100001011010010101001001001011010010100110110;
sorted_eigen_vectors[11][7] = 64'b1011111110011000001010111100011000100111111001100010110001011011;
sorted_eigen_vectors[11][8] = 64'b1011111110001101000011111110100001100010110110100110100100000010;
sorted_eigen_vectors[11][9] = 64'b0011111110011110001110011101001000001110010100101100111001100001;
sorted_eigen_vectors[11][10] = 64'b0011111110110100110000111011111111110110100010110110010111111011;
sorted_eigen_vectors[11][11] = 64'b1011111111010110111110100001101100111100011001000011010110100110;
sorted_eigen_vectors[11][12] = 64'b0011111111100111101001110110101011000101011011000010111010110100;
sorted_eigen_vectors[11][13] = 64'b1011111111100001101110011110011000011000011011001001101100010000;
sorted_eigen_vectors[11][14] = 64'b1011111110010110000001111111110110011111101100111100010111000000;
sorted_eigen_vectors[11][15] = 64'b1011111110010001011101011101110101011011000100110010101010010110;
sorted_eigen_vectors[11][16] = 64'b1011111110001100110101101101011000111010100101100000100001000111;
sorted_eigen_vectors[11][17] = 64'b1011111101110101110101001110010010000111101010111110101100011110;
sorted_eigen_vectors[11][18] = 64'b1011111110110001001110100101110110010100111100111011111101110001;
sorted_eigen_vectors[11][19] = 64'b0011111101101010010001011000110111000111111001000001011110110010;
sorted_eigen_vectors[11][20] = 64'b1011111110101001010010001100001001110100110110110001001001010011;
sorted_eigen_vectors[11][21] = 64'b0011111101111110100011011001110010000100111111100111100001000100;
sorted_eigen_vectors[11][22] = 64'b0011111110001000110101010100111000001010101001101010000001000111;
sorted_eigen_vectors[11][23] = 64'b1011111110010010001100001000001001010101001101011111001101111011;
sorted_eigen_vectors[11][24] = 64'b1011111101101011111111010111011000000100100101010001100100010010;
sorted_eigen_vectors[11][25] = 64'b0011111101110010000001010000111111101110100100001111001101011011;
sorted_eigen_vectors[11][26] = 64'b0011111101110110110001010011011010011000110000001000110010111100;
sorted_eigen_vectors[11][27] = 64'b1011111101011000011100110011100010001100011100001010100010100100;
sorted_eigen_vectors[11][28] = 64'b1011111101101111100000111110110000100110011001010111010101101000;
sorted_eigen_vectors[11][29] = 64'b0011111100010000111001110001111001010100000111010000001000100011;
sorted_eigen_vectors[11][30] = 64'b0011111011110110000100001111011000011111111101101000010000000010;
sorted_eigen_vectors[11][31] = 64'b1011111100001110111001111001011010000011000011110111000110011100;
sorted_eigen_vectors[12][0] = 64'b1011111101110100110101111100111001001100010101011100000110111001;
sorted_eigen_vectors[12][1] = 64'b1011111111000101111111001001110110110000111010000000110011101101;
sorted_eigen_vectors[12][2] = 64'b1011111111010101100111001010110101001110000101101111001000011001;
sorted_eigen_vectors[12][3] = 64'b1011111110101010000111111011110100000101011100010001100010010010;
sorted_eigen_vectors[12][4] = 64'b1011111110100001110000111110110000110000000101110100001000101010;
sorted_eigen_vectors[12][5] = 64'b0011111110100100101011011111000101001111100010010010101100100010;
sorted_eigen_vectors[12][6] = 64'b0011111110111000010101110010110011110010000110011100101011100111;
sorted_eigen_vectors[12][7] = 64'b1011111111000111010100001011000011010011110010111101111100111010;
sorted_eigen_vectors[12][8] = 64'b0011111111000101001001101001110011111010010010001110000111001100;
sorted_eigen_vectors[12][9] = 64'b1011111111001001000110000101010101110111111110100000111110101110;
sorted_eigen_vectors[12][10] = 64'b0011111110111101111000111110100100010010001000001001100101000110;
sorted_eigen_vectors[12][11] = 64'b1011111110010100010110101101000010000001010001100101010100111000;
sorted_eigen_vectors[12][12] = 64'b1011111110101101101111011101010011001110111001011010010001110110;
sorted_eigen_vectors[12][13] = 64'b1011111110001000100101100010101101101101011011110001000000100110;
sorted_eigen_vectors[12][14] = 64'b1011111110011100011010110011110000100000011110001001101000010011;
sorted_eigen_vectors[12][15] = 64'b1011111110101010100111110000010111010011000101111110001011100010;
sorted_eigen_vectors[12][16] = 64'b0011111111000011001011100010011011010100100001100011010101111110;
sorted_eigen_vectors[12][17] = 64'b1011111111011101110010101011000001001100000111001110101100010101;
sorted_eigen_vectors[12][18] = 64'b1011111111011101001001011110111001111101111001001111000001100011;
sorted_eigen_vectors[12][19] = 64'b1011111111011011000011011100010001000011000100010110010110001111;
sorted_eigen_vectors[12][20] = 64'b0011111110111010110111101101110010011111010100111111010101000001;
sorted_eigen_vectors[12][21] = 64'b1011111110100111000100100110101011111010100001100000001100011101;
sorted_eigen_vectors[12][22] = 64'b0011111110110001111110001111100110111111010000010110111011011010;
sorted_eigen_vectors[12][23] = 64'b0011111111010001111001100011111011001101001010101011100100110011;
sorted_eigen_vectors[12][24] = 64'b1011111110000010100111100001000100110011000101111001000001010110;
sorted_eigen_vectors[12][25] = 64'b1011111110000101110010110101010011000010000111111111010101100000;
sorted_eigen_vectors[12][26] = 64'b1011111101110010101101110110010011011101011010001111101000001100;
sorted_eigen_vectors[12][27] = 64'b1011111101111111010010100101011000000001100001000011000111011010;
sorted_eigen_vectors[12][28] = 64'b0011111110000000111100010110100110101111011011100100011011100111;
sorted_eigen_vectors[12][29] = 64'b1011111101100111110001011111101011100010001001011010111100000011;
sorted_eigen_vectors[12][30] = 64'b0011111101110001101101110110001000100101010100011101011011010110;
sorted_eigen_vectors[12][31] = 64'b0011111110001100100011110010011111010110100110010010000100000111;
sorted_eigen_vectors[13][0] = 64'b0011111111000000100011010001110000101101000110010111100001111110;
sorted_eigen_vectors[13][1] = 64'b0011111111000100101001010111111010111001011110000010101001100010;
sorted_eigen_vectors[13][2] = 64'b1011111110110111001111000111000110111001001101101100010011000100;
sorted_eigen_vectors[13][3] = 64'b1011111111010011001000111001101111000111011111010010000010101011;
sorted_eigen_vectors[13][4] = 64'b0011111111011111110010011110010100001000010010011011101111101000;
sorted_eigen_vectors[13][5] = 64'b0011111110010000010100100001011110110111000010001100110010010010;
sorted_eigen_vectors[13][6] = 64'b0011111110100100010111001111010000111100101011110000011001110111;
sorted_eigen_vectors[13][7] = 64'b0011111111000010001011101001010010100110011101010100001010111111;
sorted_eigen_vectors[13][8] = 64'b0011111110100111110100110001110010101111010001100110100000100010;
sorted_eigen_vectors[13][9] = 64'b0011111110101001000101110000101011001011101000001010011111010000;
sorted_eigen_vectors[13][10] = 64'b0011111110100010011100100101001101010100011010100101001011010000;
sorted_eigen_vectors[13][11] = 64'b1011111111000001001000111010111000001100010100100010000011110001;
sorted_eigen_vectors[13][12] = 64'b1011111110110001001101111111010000010011011001011001001001100100;
sorted_eigen_vectors[13][13] = 64'b0011111101110111100010000100101101111000110001100101100011000110;
sorted_eigen_vectors[13][14] = 64'b1011111111001011011000100001010110001011000101100111001101011100;
sorted_eigen_vectors[13][15] = 64'b1011111110101110110100011001011001111111001111111111000101110000;
sorted_eigen_vectors[13][16] = 64'b1011111110010010110101010111110101110001101111010001100111000101;
sorted_eigen_vectors[13][17] = 64'b1011111110001100010001010110001011100000011101010001000011111001;
sorted_eigen_vectors[13][18] = 64'b0011111101111001000000100110110001111110101110011110100001010101;
sorted_eigen_vectors[13][19] = 64'b1011111110000101101000101000101000001101111110110110001111100001;
sorted_eigen_vectors[13][20] = 64'b0011111101111110111101001010000010100111011010100001111110001110;
sorted_eigen_vectors[13][21] = 64'b0011111111000010100001101001001011100001010101000010111000110011;
sorted_eigen_vectors[13][22] = 64'b0011111110100000111101111100000110111111010000000111111100110010;
sorted_eigen_vectors[13][23] = 64'b0011111110001100100111011100100011000000010010010100101011001111;
sorted_eigen_vectors[13][24] = 64'b0011111110110100000111001110010100000111100010011010001100011010;
sorted_eigen_vectors[13][25] = 64'b0011111101110110110110000001000101000011110110111000001110100001;
sorted_eigen_vectors[13][26] = 64'b1011111101110101100000001110000000000010110101101011000101001000;
sorted_eigen_vectors[13][27] = 64'b0011111110011000111010101111110110000011010010000111001110001100;
sorted_eigen_vectors[13][28] = 64'b0011111110010011110100111101101111111000100010100001011110100001;
sorted_eigen_vectors[13][29] = 64'b0011111111100110001011101111100010000110001010000011010100111101;
sorted_eigen_vectors[13][30] = 64'b0011111110101001000000000001000110111010010011111010011110110111;
sorted_eigen_vectors[13][31] = 64'b1011111100000101100001101101110011000000010101110011011110000010;
sorted_eigen_vectors[14][0] = 64'b0011111111000001100001000110010011111110101111011011111011111000;
sorted_eigen_vectors[14][1] = 64'b0011111111000111000100101111101010010111011011001101010000000000;
sorted_eigen_vectors[14][2] = 64'b1011111110111001111111011010100010011111000100110100111110001010;
sorted_eigen_vectors[14][3] = 64'b1011111111010010111101011011000011001110110000010100011010000000;
sorted_eigen_vectors[14][4] = 64'b0011111111011110111101000011011100110110111101101110000101100110;
sorted_eigen_vectors[14][5] = 64'b0011111110100000110011001110001101111010111110000110101100010000;
sorted_eigen_vectors[14][6] = 64'b0011111110100111100001000011101011011010111000011110101110001011;
sorted_eigen_vectors[14][7] = 64'b0011111111000010110111000111100001001011000111111000001110001111;
sorted_eigen_vectors[14][8] = 64'b0011111110100111001000111101101111001010000110000000011011011100;
sorted_eigen_vectors[14][9] = 64'b0011111110100111010111000000000100000111010110110010001110011000;
sorted_eigen_vectors[14][10] = 64'b0011111110100001000100111101111111001101110111101000100111110001;
sorted_eigen_vectors[14][11] = 64'b1011111110111110110010001001011001101011100010110010111100110010;
sorted_eigen_vectors[14][12] = 64'b1011111110110000100011110010101111110110011011100000111100110010;
sorted_eigen_vectors[14][13] = 64'b0011111100111010111011010101101001011101001100101001111111100000;
sorted_eigen_vectors[14][14] = 64'b1011111111001001111111001000001111101011010011000000011111100101;
sorted_eigen_vectors[14][15] = 64'b1011111110101101010000011110100011100001110101100010100010100011;
sorted_eigen_vectors[14][16] = 64'b1011111110010100110110000011110010100000110001111101010110010110;
sorted_eigen_vectors[14][17] = 64'b1011111101010100100001011101110100111011010001011010011100101100;
sorted_eigen_vectors[14][18] = 64'b1011111101101101100101001100101111011111111110100001110001011111;
sorted_eigen_vectors[14][19] = 64'b1011111101100011110100101001101000101101110011111111111000110000;
sorted_eigen_vectors[14][20] = 64'b0011111110010100100100101011101011110101010101000000100000011111;
sorted_eigen_vectors[14][21] = 64'b0011111110111100001101011010110110111100010011001011110010100110;
sorted_eigen_vectors[14][22] = 64'b0011111110100110110010100100000111001010110111110010100011101001;
sorted_eigen_vectors[14][23] = 64'b1011111101010010011011110000001010000110101001110001101101001101;
sorted_eigen_vectors[14][24] = 64'b1011111110110101011011010001001111011010001100100110001010110101;
sorted_eigen_vectors[14][25] = 64'b0011111101100011100101010000100011101100110111011010001001000110;
sorted_eigen_vectors[14][26] = 64'b1011111110000010000000011100010110011111110011110101000011001000;
sorted_eigen_vectors[14][27] = 64'b1011111110100101101101111110101111010010110000111111000000000100;
sorted_eigen_vectors[14][28] = 64'b1011111110000000001010101110000111010111010000001011000011110100;
sorted_eigen_vectors[14][29] = 64'b1011111111100110100100000100110011000100010110100111100010001111;
sorted_eigen_vectors[14][30] = 64'b1011111110101001001100010010011011011011101000100010001100110101;
sorted_eigen_vectors[14][31] = 64'b0011111100110000011000110100001111101100010000111001110111111100;
sorted_eigen_vectors[15][0] = 64'b1011111101110010001010111001000110111100110110011001100111111100;
sorted_eigen_vectors[15][1] = 64'b1011111110110100101110011100110011100101111010001001101111010000;
sorted_eigen_vectors[15][2] = 64'b1011111110100001110111010010010000000001100011000100101101010010;
sorted_eigen_vectors[15][3] = 64'b0011111111011111011111101110001110011110110000100011111001101101;
sorted_eigen_vectors[15][4] = 64'b0011111111010011111001110001010011100110111110110101000011110001;
sorted_eigen_vectors[15][5] = 64'b1011111111010000001001010001010110100111010100100101111011101000;
sorted_eigen_vectors[15][6] = 64'b0011111110110100011101100110001010100000111010001001110000100001;
sorted_eigen_vectors[15][7] = 64'b0011111111000011011001000010001000000000000000001100010010110111;
sorted_eigen_vectors[15][8] = 64'b0011111111000000111100100101111001001001111001110001010100100000;
sorted_eigen_vectors[15][9] = 64'b1011111110000110000100111001101000100100011101111100001110110010;
sorted_eigen_vectors[15][10] = 64'b0011111110100101011011111111101011010111011010010110101010111110;
sorted_eigen_vectors[15][11] = 64'b0011111111000100111010001111010000010010101011010000101000010101;
sorted_eigen_vectors[15][12] = 64'b0011111110110000000110001100010001101110011000111011101111011110;
sorted_eigen_vectors[15][13] = 64'b1011111110011110011001111010100011001100100011100000001010100101;
sorted_eigen_vectors[15][14] = 64'b1011111110100001001000110000100001000101100011010110110001100011;
sorted_eigen_vectors[15][15] = 64'b1011111110010000001101001110000000010011011100110011011011110001;
sorted_eigen_vectors[15][16] = 64'b0011111110110000001001111001110010111110010001011011000100010010;
sorted_eigen_vectors[15][17] = 64'b1011111110010100010101001010100011010110010101110110110010011110;
sorted_eigen_vectors[15][18] = 64'b0011111101101000100100111110000100011001001011010000111101110011;
sorted_eigen_vectors[15][19] = 64'b1011111110010100000011101011100110000011101110000011111100010010;
sorted_eigen_vectors[15][20] = 64'b1011111110110100011101110010011101101010001010011001110100000011;
sorted_eigen_vectors[15][21] = 64'b0011111110011000010100110101100000111001001011010110110101101101;
sorted_eigen_vectors[15][22] = 64'b1011111110100010100011010100101110000000101110110110011010011000;
sorted_eigen_vectors[15][23] = 64'b0011111110011011111001000100111110100001100010110011110000100100;
sorted_eigen_vectors[15][24] = 64'b0011111110111010000101111111011010101111110111100011111111101110;
sorted_eigen_vectors[15][25] = 64'b0011111110110101111000010011011010100010011010011110101100001111;
sorted_eigen_vectors[15][26] = 64'b1011111111000111010101010010001100100010101001011000100111111011;
sorted_eigen_vectors[15][27] = 64'b0011111111100101000000001000110001010111000100110110110111101011;
sorted_eigen_vectors[15][28] = 64'b0011111110110110011101110000001101111001010100000111110011001111;
sorted_eigen_vectors[15][29] = 64'b1011111110101011011011111111001000010101010000110101000010011111;
sorted_eigen_vectors[15][30] = 64'b0011111110100111000011001001111010101000101000010000010000001111;
sorted_eigen_vectors[15][31] = 64'b0011111100010000101111110111110001111101101100010100110010011001;
sorted_eigen_vectors[16][0] = 64'b1011111110001010011100000100111011100011001011111111101100011000;
sorted_eigen_vectors[16][1] = 64'b1011111110110010011011101010011100001111000011001101010010101011;
sorted_eigen_vectors[16][2] = 64'b1011111110100110000110111000110110011110011010011101101001010000;
sorted_eigen_vectors[16][3] = 64'b0011111111011111100010110010000010010110101100011110101000111011;
sorted_eigen_vectors[16][4] = 64'b0011111111010011010110010101010100011100011110100000011001010100;
sorted_eigen_vectors[16][5] = 64'b1011111111001110110101110110011010110001110011101010010100110010;
sorted_eigen_vectors[16][6] = 64'b0011111110110110010101101100110011011000000001011000000000001110;
sorted_eigen_vectors[16][7] = 64'b0011111111000101001101111000110110001101101010000100001111010010;
sorted_eigen_vectors[16][8] = 64'b0011111111000010101001100111011000011110010001111000010000101100;
sorted_eigen_vectors[16][9] = 64'b1011111110001110010010001001111100001110001001011011110001010001;
sorted_eigen_vectors[16][10] = 64'b0011111110101010111100101000001110011011010101110100110000100000;
sorted_eigen_vectors[16][11] = 64'b0011111111000110010110000111111010001101000110111110100010000010;
sorted_eigen_vectors[16][12] = 64'b0011111110110100100110100110111000101001100100011011000010100000;
sorted_eigen_vectors[16][13] = 64'b1011111110010010000001011100100000110110100011110100011011010011;
sorted_eigen_vectors[16][14] = 64'b1011111110010100110001001000110110001111011111100011010100111011;
sorted_eigen_vectors[16][15] = 64'b1011111110001000010101110111100011010101100111000000011000011001;
sorted_eigen_vectors[16][16] = 64'b0011111110110010111100101101010110111101100101101000101001000011;
sorted_eigen_vectors[16][17] = 64'b0011111110100011111110011101011110000001111011111000100111100101;
sorted_eigen_vectors[16][18] = 64'b1011111110000101111000110101110001101000101111110111011111011100;
sorted_eigen_vectors[16][19] = 64'b1011111101110110011001011101101111100001110100101011011110101111;
sorted_eigen_vectors[16][20] = 64'b0011111110110101001101111001000010001011000100001110010100111100;
sorted_eigen_vectors[16][21] = 64'b1011111110001111001100100100010101011111101000101011011100101000;
sorted_eigen_vectors[16][22] = 64'b1011111101110110001101011100011110010000101011010011010010001100;
sorted_eigen_vectors[16][23] = 64'b1011111100010100011010101010011111101010111010110101110111110000;
sorted_eigen_vectors[16][24] = 64'b1011111111000000000110100010111110000110110110011100101100001111;
sorted_eigen_vectors[16][25] = 64'b1011111110101001011110000001011001110111110000101111001010100010;
sorted_eigen_vectors[16][26] = 64'b0011111111000101110100111000010111110100101011101100011111110011;
sorted_eigen_vectors[16][27] = 64'b1011111111100100111100111100011100010011011110111000101111010000;
sorted_eigen_vectors[16][28] = 64'b1011111110110111001111011000000111100000001010001101111100000110;
sorted_eigen_vectors[16][29] = 64'b0011111110101001001000111101110001000110100010010000010001100000;
sorted_eigen_vectors[16][30] = 64'b1011111110101000011001110101111000111011011001100101010100111100;
sorted_eigen_vectors[16][31] = 64'b1011111100110100011000010001010011100010010011110001111010111101;
sorted_eigen_vectors[17][0] = 64'b1011111111011101111010000001100000001111000101110101110100101001;
sorted_eigen_vectors[17][1] = 64'b0011111110100111100100011100001101100010011001010010010001101101;
sorted_eigen_vectors[17][2] = 64'b1011111101111110111110110111100111101000100110010001011111111111;
sorted_eigen_vectors[17][3] = 64'b1011111110110110011110010110000100100101000110001110001011000001;
sorted_eigen_vectors[17][4] = 64'b0011111110111110000001110111100000111110011100111010101000011011;
sorted_eigen_vectors[17][5] = 64'b1011111110001111000011010100000100000000010000101000100101011011;
sorted_eigen_vectors[17][6] = 64'b1011111110100011011010010010011110010011001011111111001110000110;
sorted_eigen_vectors[17][7] = 64'b1011111110101110001010100000001001010100111110110011110110001101;
sorted_eigen_vectors[17][8] = 64'b1011111110100100110000000101000101110010101100100101011010110011;
sorted_eigen_vectors[17][9] = 64'b1011111101110010110111110101010110010110111011011001111110100001;
sorted_eigen_vectors[17][10] = 64'b0011111110010110001010101010100000101000010111111001000100001001;
sorted_eigen_vectors[17][11] = 64'b0011111110110011111011111001001001010010111110000010011111010010;
sorted_eigen_vectors[17][12] = 64'b0011111101110000000111100111110011100001010001000111101110001111;
sorted_eigen_vectors[17][13] = 64'b1011111110101000100101111101001100001000000101011111111001000011;
sorted_eigen_vectors[17][14] = 64'b0011111110101011101111010110000111111011000000000000110011010011;
sorted_eigen_vectors[17][15] = 64'b0011111110010001001100011000000100001011110111110110101110110000;
sorted_eigen_vectors[17][16] = 64'b1011111110100010111000100010000011101000100111011010001011101011;
sorted_eigen_vectors[17][17] = 64'b1011111110011011111100100000010111001000000100111111001011111011;
sorted_eigen_vectors[17][18] = 64'b0011111110100001111111011010001101111001101010111100001000010000;
sorted_eigen_vectors[17][19] = 64'b1011111101111100110010010110011101001010000010100011010110100100;
sorted_eigen_vectors[17][20] = 64'b0011111110011001100101001011011001011011000100100001000110011011;
sorted_eigen_vectors[17][21] = 64'b0011111110001011110101101000000100100001111101111110111010111001;
sorted_eigen_vectors[17][22] = 64'b1011111110100111110110101010000111101101010111010100010111100101;
sorted_eigen_vectors[17][23] = 64'b0011111110100011011000001001111000100011011001111000010000001110;
sorted_eigen_vectors[17][24] = 64'b1011111110101110011010000001000000000001010010101100010111101101;
sorted_eigen_vectors[17][25] = 64'b0011111111011100111000110010010101000011010110111001100011011110;
sorted_eigen_vectors[17][26] = 64'b1011111110100010101000101010000001010010000111000101110101010101;
sorted_eigen_vectors[17][27] = 64'b1011111110110111100100110011101001010000000001111000010101011110;
sorted_eigen_vectors[17][28] = 64'b1011111110101001000111010101001011011101111100001110010001101101;
sorted_eigen_vectors[17][29] = 64'b1011111110100101101101011100000011100010000001000010001000011010;
sorted_eigen_vectors[17][30] = 64'b0011111111100110110110101001000011111101000010111011110000000101;
sorted_eigen_vectors[17][31] = 64'b0011111101010000010100111010001010100111011010110001011110100010;
sorted_eigen_vectors[18][0] = 64'b1011111111011101101111000000011011001011011001011110011010000111;
sorted_eigen_vectors[18][1] = 64'b0011111110100110111110100000011100000011000111101110001101010100;
sorted_eigen_vectors[18][2] = 64'b1011111101111101010100100110011011011000110001100001001110101010;
sorted_eigen_vectors[18][3] = 64'b1011111110110111100110101001101011110001101011010001100010100011;
sorted_eigen_vectors[18][4] = 64'b0011111110111110000011101010000101111001101100000100100101010111;
sorted_eigen_vectors[18][5] = 64'b1011111110010000010001100111000111000000101010110001101010100010;
sorted_eigen_vectors[18][6] = 64'b1011111110100100100100110011001010011011000001001011111101010000;
sorted_eigen_vectors[18][7] = 64'b1011111110110000101010110100010110000110110101011111001111110011;
sorted_eigen_vectors[18][8] = 64'b1011111110100101100101111000001011010010111111101000000000001001;
sorted_eigen_vectors[18][9] = 64'b1011111101111110001010110001100100111101000001001110100101011100;
sorted_eigen_vectors[18][10] = 64'b0011111110010100001111100011001011001101110010100000100010100110;
sorted_eigen_vectors[18][11] = 64'b0011111110110101000111110111000110010101111110011101111111110100;
sorted_eigen_vectors[18][12] = 64'b0011111101110001110000101100101100100011011011001010100110010100;
sorted_eigen_vectors[18][13] = 64'b1011111110101001011111001010011111011110100001011100011010000011;
sorted_eigen_vectors[18][14] = 64'b0011111110101011100110010000010011110011000110100110011101110100;
sorted_eigen_vectors[18][15] = 64'b0011111110010000110000000101010010011010110001100010111010111101;
sorted_eigen_vectors[18][16] = 64'b1011111110100011100010000011010011000100000011001011101000011100;
sorted_eigen_vectors[18][17] = 64'b1011111110011011111111010000000000001010001001100011111010111011;
sorted_eigen_vectors[18][18] = 64'b0011111110011010011001111100100100010000100100110110010101010111;
sorted_eigen_vectors[18][19] = 64'b1011111101111000011110111100001110011110110001010101101010000011;
sorted_eigen_vectors[18][20] = 64'b0011111110010111100101110111111011100101100010100000111001010010;
sorted_eigen_vectors[18][21] = 64'b0011111110011011010011101001001011101100101010010101111111011111;
sorted_eigen_vectors[18][22] = 64'b1011111110101100100010111011100010110110000101011101101111110101;
sorted_eigen_vectors[18][23] = 64'b0011111110101011001101010100011110111010110000110110101010100101;
sorted_eigen_vectors[18][24] = 64'b1011111110100101101111101010011000000010000010000010101010111101;
sorted_eigen_vectors[18][25] = 64'b0011111111011111101110110010110110111011100000100010100010110010;
sorted_eigen_vectors[18][26] = 64'b1011111110000001001000000000010011100000001001001001100100100100;
sorted_eigen_vectors[18][27] = 64'b0011111110000001101101100001010110010110101101000100000001001111;
sorted_eigen_vectors[18][28] = 64'b1011111110001111100110110010011110111001111100001100000011101000;
sorted_eigen_vectors[18][29] = 64'b0011111110101000100110111001010110100000000011010011010001111101;
sorted_eigen_vectors[18][30] = 64'b1011111111100110001000110100000100100110010001100111010001101010;
sorted_eigen_vectors[18][31] = 64'b1011111101011000010001100011100100011001000000010100111100110000;
sorted_eigen_vectors[19][0] = 64'b1011111110011101001000001010000111000100000010010100101110010100;
sorted_eigen_vectors[19][1] = 64'b0011111111001111100100110011010111001000000111110100010011000100;
sorted_eigen_vectors[19][2] = 64'b1011111111001001000001010000111010100111000111001101100011110101;
sorted_eigen_vectors[19][3] = 64'b0011111111000100011010001010011111101000010000111011010100111000;
sorted_eigen_vectors[19][4] = 64'b1011111110110011011011110010101101110011001010101000110001000000;
sorted_eigen_vectors[19][5] = 64'b0011111111011101000000111010011000000100001110111100100111110001;
sorted_eigen_vectors[19][6] = 64'b0011111111000100000001010110111100001000001010001001100100010110;
sorted_eigen_vectors[19][7] = 64'b0011111111001110000101010011001010011110110100001011001111000100;
sorted_eigen_vectors[19][8] = 64'b1011111110110111100101000011011111101101010100001101011011100000;
sorted_eigen_vectors[19][9] = 64'b0011111110101111011100000100111000000011101101101110011101010011;
sorted_eigen_vectors[19][10] = 64'b0011111111000000010001100111011100011000111110100110010110000010;
sorted_eigen_vectors[19][11] = 64'b0011111110110101111001111100111110101000000000000110101101101001;
sorted_eigen_vectors[19][12] = 64'b1011111110101011001101001110111101001010001011100000111101001101;
sorted_eigen_vectors[19][13] = 64'b1011111110111101000110101110010100001010011010010011010000111111;
sorted_eigen_vectors[19][14] = 64'b0011111110110010111010010001110001111000011001100111100111010110;
sorted_eigen_vectors[19][15] = 64'b0011111110011000100101001110111010101110001100101100011010010011;
sorted_eigen_vectors[19][16] = 64'b0011111110111010011000110100100010001111100010101000110000000110;
sorted_eigen_vectors[19][17] = 64'b0011111110010101110100000010101001101110110100001111001111010010;
sorted_eigen_vectors[19][18] = 64'b0011111110100000101110100010110101000110010101111101111001110001;
sorted_eigen_vectors[19][19] = 64'b1011111110010001110110110010110011001011110111011011111000100111;
sorted_eigen_vectors[19][20] = 64'b0011111110101011010101100001111101100101000010011001111000110011;
sorted_eigen_vectors[19][21] = 64'b1011111110011010010001011011110001110011001110111011101100110010;
sorted_eigen_vectors[19][22] = 64'b0011111110100010000001001110100101111001011101001100110111111011;
sorted_eigen_vectors[19][23] = 64'b1011111110100000101110011111011010110010100001100000000110001110;
sorted_eigen_vectors[19][24] = 64'b1011111111100110000011111100111000101001111100001100000100001100;
sorted_eigen_vectors[19][25] = 64'b1011111110100111001101010100001110001100001010010111010000101100;
sorted_eigen_vectors[19][26] = 64'b1011111110101110011010011000101011110011111011110110010010111110;
sorted_eigen_vectors[19][27] = 64'b0011111111000000100101010101100100000011101011000110100011101011;
sorted_eigen_vectors[19][28] = 64'b0011111110101000111100100001010000010111010011011010001011110111;
sorted_eigen_vectors[19][29] = 64'b0011111110110110101101101111010001001100001100111100101000101111;
sorted_eigen_vectors[19][30] = 64'b0011111101011110110011110000000000101110011000111011101000001010;
sorted_eigen_vectors[19][31] = 64'b0011111101000010010111100110101101101011011010100111110010111000;
sorted_eigen_vectors[20][0] = 64'b0011111110010111110110110001010110111111001001000011110110101100;
sorted_eigen_vectors[20][1] = 64'b1011111111001110101100110101010011111111111100001100001001000010;
sorted_eigen_vectors[20][2] = 64'b0011111111001000100110101000100111011111000010010100001000111011;
sorted_eigen_vectors[20][3] = 64'b1011111111000100101011110110100100111010111101011110001010110101;
sorted_eigen_vectors[20][4] = 64'b0011111110101010101101000010111100110000001101100100110001001111;
sorted_eigen_vectors[20][5] = 64'b1011111111011100110111101111011100110100110011001000101111110111;
sorted_eigen_vectors[20][6] = 64'b1011111111000100001011111010110111111000010011011111001010001000;
sorted_eigen_vectors[20][7] = 64'b1011111111001110000011111111100111001101111110111011100011100001;
sorted_eigen_vectors[20][8] = 64'b0011111110111010010000010010111100011000001111000101001000100110;
sorted_eigen_vectors[20][9] = 64'b1011111110110000000110000110101111000100001001011101010100000100;
sorted_eigen_vectors[20][10] = 64'b1011111111000000101110010110110111110101101101001101100010001010;
sorted_eigen_vectors[20][11] = 64'b1011111110110110110011011110000111110001110000001111111100110101;
sorted_eigen_vectors[20][12] = 64'b0011111110101011110111011110000100110000001100101111100111010011;
sorted_eigen_vectors[20][13] = 64'b0011111111000001000110101001110011001111100111101000101101111011;
sorted_eigen_vectors[20][14] = 64'b1011111110111001001010001001011010100000100110011100010101111011;
sorted_eigen_vectors[20][15] = 64'b1011111110100011001011001000101101110100111001111001101010101000;
sorted_eigen_vectors[20][16] = 64'b1011111111000010010111000001110011111010011110100111001000011100;
sorted_eigen_vectors[20][17] = 64'b0011111101110000000000101001111110001011011001100011111011011101;
sorted_eigen_vectors[20][18] = 64'b1011111110110101011110000100100101001010010111101100011111000011;
sorted_eigen_vectors[20][19] = 64'b0011111110101100010001100101000000001110010001010010110100101101;
sorted_eigen_vectors[20][20] = 64'b1011111110100000011101000011011011100011000111111000100010110010;
sorted_eigen_vectors[20][21] = 64'b1011111101000000001000110100100111010010001100110111010010110101;
sorted_eigen_vectors[20][22] = 64'b0011111110111011110000111010000111010011110110010110111001101110;
sorted_eigen_vectors[20][23] = 64'b1011111110100001110010011101111001011000100010110101010101001010;
sorted_eigen_vectors[20][24] = 64'b1011111111100101101000011001000001101110111110100101111110100101;
sorted_eigen_vectors[20][25] = 64'b1011111110101011000011100010111110110111000011001000010110010111;
sorted_eigen_vectors[20][26] = 64'b1011111110101010000111001011100100101111001110111110010110100110;
sorted_eigen_vectors[20][27] = 64'b0011111110111010001010100001111010101000001110001000001101000011;
sorted_eigen_vectors[20][28] = 64'b0011111101111000011000010010110000110000111101101001110100000000;
sorted_eigen_vectors[20][29] = 64'b0011111110101111011011001110111011000101010111001010110001101101;
sorted_eigen_vectors[20][30] = 64'b0011111101100011011101100001011010100110011100110000110100011110;
sorted_eigen_vectors[20][31] = 64'b0011111100110001001101001100101101111100111011101101011000010111;
sorted_eigen_vectors[21][0] = 64'b1011111110110001011010111010000111001111010000010010111001101011;
sorted_eigen_vectors[21][1] = 64'b0011111110001110101111010111001111101110000100100110000110011010;
sorted_eigen_vectors[21][2] = 64'b0011111110000010111100100010110011110111100010000001111001011101;
sorted_eigen_vectors[21][3] = 64'b0011111110111101100011010101100101010101000001110100010100101101;
sorted_eigen_vectors[21][4] = 64'b1011111111000110010001100100110100101000010101000000001110100101;
sorted_eigen_vectors[21][5] = 64'b1011111110100000001001101110101001101110110100101010001001110000;
sorted_eigen_vectors[21][6] = 64'b1011111101111000001000001111101001111101000110010100010100001100;
sorted_eigen_vectors[21][7] = 64'b1011111110111000010000110101000000101111011010001110101010101001;
sorted_eigen_vectors[21][8] = 64'b1011111110110110100101001000001111110110101111011101010110000001;
sorted_eigen_vectors[21][9] = 64'b1011111110100101011100011100000111010111111000010111001101110000;
sorted_eigen_vectors[21][10] = 64'b1011111110100001011110000100100110010000000011100001110001101011;
sorted_eigen_vectors[21][11] = 64'b0011111110111100110111101111010000001111010100111100001111101100;
sorted_eigen_vectors[21][12] = 64'b1011111111010101111101001000011011001111111011101100100010011100;
sorted_eigen_vectors[21][13] = 64'b1011111111011111010001100101001010111000111011111000001100110000;
sorted_eigen_vectors[21][14] = 64'b1011111111100110101101001011110100000001111011011101010001000011;
sorted_eigen_vectors[21][15] = 64'b1011111110111110111010010001111101000011010001011110100001101001;
sorted_eigen_vectors[21][16] = 64'b1011111110111111100000010110110010101111101110000000010000011010;
sorted_eigen_vectors[21][17] = 64'b0011111110110010100011101011110101011010110001001100100011101100;
sorted_eigen_vectors[21][18] = 64'b1011111110110001100000011001001110101001001001010010101011000110;
sorted_eigen_vectors[21][19] = 64'b0011111110101101101011011010001011100000111001100100000001010111;
sorted_eigen_vectors[21][20] = 64'b1011111110110000110101100111110111000011011100001111000111100001;
sorted_eigen_vectors[21][21] = 64'b1011111110111000011010101110010110010011001000100010100101000110;
sorted_eigen_vectors[21][22] = 64'b1011111110100000010011111101011011101101001111000011111010100100;
sorted_eigen_vectors[21][23] = 64'b0011111101101011101101001001010010101110101101000011010110000110;
sorted_eigen_vectors[21][24] = 64'b0011111110000111011101101000011001111000011001001110110001101001;
sorted_eigen_vectors[21][25] = 64'b1011111101011011010000000011101010011011111110010010011001101111;
sorted_eigen_vectors[21][26] = 64'b0011111110000011111000010101100100011111000111000110100110001011;
sorted_eigen_vectors[21][27] = 64'b1011111110010011001001011011010011110111110011110011100100110111;
sorted_eigen_vectors[21][28] = 64'b0011111101110001000010000110110100111000101111110000010011100110;
sorted_eigen_vectors[21][29] = 64'b0011111100100111111100011111000010001111011010010011011101100011;
sorted_eigen_vectors[21][30] = 64'b0011111100110101001010010100110100000110101001100001010111100111;
sorted_eigen_vectors[21][31] = 64'b1011111100110011001011011000000010011011010011010001101001001100;
sorted_eigen_vectors[22][0] = 64'b0011111111001010010011011011110011010101100111011001111001000000;
sorted_eigen_vectors[22][1] = 64'b1011111110000001000111011011110111101111011000001101100100111000;
sorted_eigen_vectors[22][2] = 64'b0011111101100111100100011001101001011000110100011110011101011100;
sorted_eigen_vectors[22][3] = 64'b1011111111001000001011011101101101000110010110111100000011111111;
sorted_eigen_vectors[22][4] = 64'b0011111111010010010110100001000110100111111011100000111101101010;
sorted_eigen_vectors[22][5] = 64'b1011111110011011101000100111100111011110110100110100100111101111;
sorted_eigen_vectors[22][6] = 64'b1011111110111011011111101001101101111011001000010110010111010001;
sorted_eigen_vectors[22][7] = 64'b1011111111001100010001110011011000001011110110011111100010010110;
sorted_eigen_vectors[22][8] = 64'b1011111111000101001110011101011000001111011111011010100010010001;
sorted_eigen_vectors[22][9] = 64'b1011111110010011110100010100001110010010100011101110100101010101;
sorted_eigen_vectors[22][10] = 64'b0011111110110101001101000100100111000111010011011111101110001101;
sorted_eigen_vectors[22][11] = 64'b0011111111010001100111000001011001111001001000101010101111010001;
sorted_eigen_vectors[22][12] = 64'b1011111110100101111110110101010010010101001000101110001010011011;
sorted_eigen_vectors[22][13] = 64'b1011111111001100000010111101110110011101000100100010110010100100;
sorted_eigen_vectors[22][14] = 64'b0011111111001010101010101011111011001000001101011110011011111111;
sorted_eigen_vectors[22][15] = 64'b0011111110111100100010000111111001111001001110011110110101110000;
sorted_eigen_vectors[22][16] = 64'b0011111111010001010100011000010011101010101110100110101011111110;
sorted_eigen_vectors[22][17] = 64'b0011111111000100100010100111010011100011100011110011100000001100;
sorted_eigen_vectors[22][18] = 64'b1011111110111001000000100110110011000101100011010010110010110001;
sorted_eigen_vectors[22][19] = 64'b0011111110011110100001101000000011111000111001111011100110110000;
sorted_eigen_vectors[22][20] = 64'b1011111110111101001110101100010111001100111001001000001111101011;
sorted_eigen_vectors[22][21] = 64'b1011111111100011111010100101100100011111101110110110110100111101;
sorted_eigen_vectors[22][22] = 64'b1011111111001001010110001000100011001001100010111110100001000010;
sorted_eigen_vectors[22][23] = 64'b1011111101110000001010010110001001101010010111001100001111000110;
sorted_eigen_vectors[22][24] = 64'b1011111110011010010011001110101011000111001111100100000101111010;
sorted_eigen_vectors[22][25] = 64'b1011111110000100111010010101011111110000000001101110000011000100;
sorted_eigen_vectors[22][26] = 64'b0011111110110001100111001000111111000000010011100001101001001000;
sorted_eigen_vectors[22][27] = 64'b0011111110100101000001101000000111101010111101101011011101011010;
sorted_eigen_vectors[22][28] = 64'b1011111110110011111011011000011001100111100010010000110101111100;
sorted_eigen_vectors[22][29] = 64'b0011111110010010111111101110010100000010101001011111001110110101;
sorted_eigen_vectors[22][30] = 64'b0011111101100100000011100010000001010011001100000111100000001100;
sorted_eigen_vectors[22][31] = 64'b1011111101001000100000100111000101001000100110011000011101000111;
sorted_eigen_vectors[23][0] = 64'b0011111110101010011001010001000100110010110000010100101111100110;
sorted_eigen_vectors[23][1] = 64'b0011111111011001110100010101011001111000011110010111101001111000;
sorted_eigen_vectors[23][2] = 64'b1011111111001010000001101001010000001111110010101110111111111011;
sorted_eigen_vectors[23][3] = 64'b0011111110101000100101011000011100011101010111101111000100010000;
sorted_eigen_vectors[23][4] = 64'b1011111110010101110100100010111011011100101010100011110001111000;
sorted_eigen_vectors[23][5] = 64'b1011111110110101001011110101100010010110011111001001011010000111;
sorted_eigen_vectors[23][6] = 64'b1011111110010001110100110111010111110110010001001000111010010011;
sorted_eigen_vectors[23][7] = 64'b1011111110111000001110101000000100100100110101101010101111000000;
sorted_eigen_vectors[23][8] = 64'b0011111110110001111010101011111100001001001000101000000111101011;
sorted_eigen_vectors[23][9] = 64'b1011111111000001001100001100010101111001100110101010011011110100;
sorted_eigen_vectors[23][10] = 64'b1011111111001001001010101010111101110011000010000100010100010100;
sorted_eigen_vectors[23][11] = 64'b0011111110111011111110101111000101000111111000010001011000000111;
sorted_eigen_vectors[23][12] = 64'b0011111110111001000110001000110111010001100101011000111010011001;
sorted_eigen_vectors[23][13] = 64'b0011111110100110110101010110100000101000011110111111011100001111;
sorted_eigen_vectors[23][14] = 64'b0011111110110101001000011111001001110011111010011010100000101001;
sorted_eigen_vectors[23][15] = 64'b0011111110010010011000000001111000100100100010101111000111011010;
sorted_eigen_vectors[23][16] = 64'b1011111111001110010100010011010110110011010000111101011111000001;
sorted_eigen_vectors[23][17] = 64'b0011111110100011110110111000010010001111100011010100100100001111;
sorted_eigen_vectors[23][18] = 64'b1011111111001000010101011011010011101111110101011110111001101001;
sorted_eigen_vectors[23][19] = 64'b0011111110111110100111001000110001001101101111101010110110001101;
sorted_eigen_vectors[23][20] = 64'b1011111111000111100011000011110101110000110001111100000010010000;
sorted_eigen_vectors[23][21] = 64'b1011111111000110111110111000110011110100111000111011111001001100;
sorted_eigen_vectors[23][22] = 64'b0011111111001111000100111111010000111101000111000011000101010011;
sorted_eigen_vectors[23][23] = 64'b1011111110011011101011111110100001101010110111011100010001100100;
sorted_eigen_vectors[23][24] = 64'b0011111110110000011110001000100111101100110100111111100111110111;
sorted_eigen_vectors[23][25] = 64'b0011111110100111111101001101001110000100000001011100011011101100;
sorted_eigen_vectors[23][26] = 64'b1011111111010111011011011000110011110100100001101001110111100001;
sorted_eigen_vectors[23][27] = 64'b1011111111001000000000100111100000101011100100001010010111101110;
sorted_eigen_vectors[23][28] = 64'b0011111111100000101101011100011011000111100011001111000110010011;
sorted_eigen_vectors[23][29] = 64'b0011111110000010001101111111001010111000101100010001011000010101;
sorted_eigen_vectors[23][30] = 64'b1011111101111010000001101000110011101000101100011101100001001001;
sorted_eigen_vectors[23][31] = 64'b0011111100101010101111010101000011100011110110110111001011001111;
sorted_eigen_vectors[24][0] = 64'b1011111110010000101011100011001000001010111101011111100100100101;
sorted_eigen_vectors[24][1] = 64'b0011111111011010011100101001100100110000010110010011101011100001;
sorted_eigen_vectors[24][2] = 64'b1011111111001010101011011010010101100001101110011000101000011001;
sorted_eigen_vectors[24][3] = 64'b0011111110110001101011111101010111000111001100111100101111011110;
sorted_eigen_vectors[24][4] = 64'b1011111110101100100011001110111001101001101100111111011010010011;
sorted_eigen_vectors[24][5] = 64'b1011111110110001110100111000111001111111110001100101011110010001;
sorted_eigen_vectors[24][6] = 64'b0011111110010101100011110110001111111001000100010100110000010001;
sorted_eigen_vectors[24][7] = 64'b1011111110001010011000110010011001111011010111101101101001100101;
sorted_eigen_vectors[24][8] = 64'b0011111110111101000110001101110111110010111001011001011011100010;
sorted_eigen_vectors[24][9] = 64'b1011111110111110010110010110010000111111001110000011110010001100;
sorted_eigen_vectors[24][10] = 64'b1011111111001001011110010110010001101110001100000101100101110110;
sorted_eigen_vectors[24][11] = 64'b0011111110011010000111101010000101001000101000001111001001010010;
sorted_eigen_vectors[24][12] = 64'b0011111110111000111101000001010001011100110110111101111011101010;
sorted_eigen_vectors[24][13] = 64'b0011111110111000101111011100110011101000101100010000101100100111;
sorted_eigen_vectors[24][14] = 64'b0011111110010110001100110100000011010000110000110011111000111111;
sorted_eigen_vectors[24][15] = 64'b1011111101111111101011010011100111100101110110111111010011001110;
sorted_eigen_vectors[24][16] = 64'b1011111111010011110111101001100011001101001101010110010111110001;
sorted_eigen_vectors[24][17] = 64'b1011111110100001101001001111101011011000111010110101101101111111;
sorted_eigen_vectors[24][18] = 64'b1011111111000000100101100011010111001000011111010110011111101110;
sorted_eigen_vectors[24][19] = 64'b0011111110110011101100000110111101011100101111110110011111000100;
sorted_eigen_vectors[24][20] = 64'b1011111110111100001100001011111110000001110011101000000100001010;
sorted_eigen_vectors[24][21] = 64'b1011111111000001101111111010011010011000100011010011100010111110;
sorted_eigen_vectors[24][22] = 64'b0011111110111100101011001011010011111110100111110010101101010110;
sorted_eigen_vectors[24][23] = 64'b1011111101110010101110101111101000111000100001000111101010100110;
sorted_eigen_vectors[24][24] = 64'b0011111110001001010110100100001110100110001110111111110001110011;
sorted_eigen_vectors[24][25] = 64'b1011111110000101110110010000001010101111111101010111101011011100;
sorted_eigen_vectors[24][26] = 64'b0011111111011001100001000111010011101110011000100101001111110111;
sorted_eigen_vectors[24][27] = 64'b0011111111000111010111001011111101000101111001001001011111101001;
sorted_eigen_vectors[24][28] = 64'b1011111111100010010110000010011111010000100010000010001111000101;
sorted_eigen_vectors[24][29] = 64'b0011111110001000111100000110100110010000110011110110100111101110;
sorted_eigen_vectors[24][30] = 64'b0011111101111100100001011101000111101101101000110110011100000101;
sorted_eigen_vectors[24][31] = 64'b1011111101011100010011011111011101000000011110111111001010010011;
sorted_eigen_vectors[25][0] = 64'b0011111101010100100000110000101100011000011100010010000110110110;
sorted_eigen_vectors[25][1] = 64'b1011111111010101100001101010011110011011000100001010111011100101;
sorted_eigen_vectors[25][2] = 64'b0011111111000111011011111000110001011110001100000101100101100010;
sorted_eigen_vectors[25][3] = 64'b1011111110111111110001111010111001100011100101000110001111011011;
sorted_eigen_vectors[25][4] = 64'b0011111110100110001101000000100101010111010100001011110110000011;
sorted_eigen_vectors[25][5] = 64'b0011111111000001110011000001000010110001011000111100011010110101;
sorted_eigen_vectors[25][6] = 64'b0011111111000011001100001110111001100110111011010000100111011000;
sorted_eigen_vectors[25][7] = 64'b0011111111001101101101111001010010001010100000100011010110000100;
sorted_eigen_vectors[25][8] = 64'b0011111110100010001100010110001001101000111011011000010100010000;
sorted_eigen_vectors[25][9] = 64'b1011111110101100000110010010011100101000001010101001110000000111;
sorted_eigen_vectors[25][10] = 64'b1011111110011101111001100011010100100100010100110101010000100010;
sorted_eigen_vectors[25][11] = 64'b0011111111000111101111110011001111011011111010010110100011001010;
sorted_eigen_vectors[25][12] = 64'b1011111110101110101001110101011111111100001111110011110000010001;
sorted_eigen_vectors[25][13] = 64'b1011111111000101001110001001101001000101010011001000111110110100;
sorted_eigen_vectors[25][14] = 64'b0011111110111001010011001001000101010110000101011000110000111011;
sorted_eigen_vectors[25][15] = 64'b0011111110100011111010000011000100000100111011000110001011100000;
sorted_eigen_vectors[25][16] = 64'b1011111110011111110110101110011100100010011101010001100010011101;
sorted_eigen_vectors[25][17] = 64'b0011111110111000100011101111001011001001000011110110000110010110;
sorted_eigen_vectors[25][18] = 64'b1011111110110101000010110100110111100100101100111011010010001111;
sorted_eigen_vectors[25][19] = 64'b0011111110001100101111001111110011000011101010101010011110110010;
sorted_eigen_vectors[25][20] = 64'b1011111110110010011111011011100011111111000111010011111000100011;
sorted_eigen_vectors[25][21] = 64'b1011111110110001111111000101111111100001011100000101000010111101;
sorted_eigen_vectors[25][22] = 64'b0011111111101000101100111000000000101101011110011111001100101100;
sorted_eigen_vectors[25][23] = 64'b1011111110110000001010000101010011010010001111100000011010100110;
sorted_eigen_vectors[25][24] = 64'b0011111110110001111111110001111101101110011001011101011110100010;
sorted_eigen_vectors[25][25] = 64'b0011111110111011111101000111001101011010111011111101000001100001;
sorted_eigen_vectors[25][26] = 64'b0011111110111011011010101011010001111001101011010011110100011101;
sorted_eigen_vectors[25][27] = 64'b0011111110011111001010111111111010110101111100001010101010111110;
sorted_eigen_vectors[25][28] = 64'b1011111110100111010100000101101011011111010111111000110111101110;
sorted_eigen_vectors[25][29] = 64'b0011111100100100110111010010011011110111110110001101111100001101;
sorted_eigen_vectors[25][30] = 64'b0011111101100001010001110100001011111010001010110101110100100000;
sorted_eigen_vectors[25][31] = 64'b1011111101001111100110110001000101001001101111100000110010100111;
sorted_eigen_vectors[26][0] = 64'b1011111110110001100010001100011110010001101110111001011000100010;
sorted_eigen_vectors[26][1] = 64'b1011111111001011100010011110101000000001110100011010010000110100;
sorted_eigen_vectors[26][2] = 64'b0011111111000010011011000011011001001001010100000000100100000011;
sorted_eigen_vectors[26][3] = 64'b1011111110111001001010011000000001111011011100101001011110000111;
sorted_eigen_vectors[26][4] = 64'b0011111110001111001111100100011011000101010110111001001100011100;
sorted_eigen_vectors[26][5] = 64'b0011111110111000100111001001000001110001111111011001111000010010;
sorted_eigen_vectors[26][6] = 64'b0011111111001011001110110001011011111000101011100110111110110111;
sorted_eigen_vectors[26][7] = 64'b0011111111011010010011100000011100010001001100100001111000000111;
sorted_eigen_vectors[26][8] = 64'b0011111111001000100010010101111101011101011110010111011011100100;
sorted_eigen_vectors[26][9] = 64'b1011111110110001111011010001111101000101010101100111101010011100;
sorted_eigen_vectors[26][10] = 64'b1011111111000101100110000000111001000111111101011010010100111010;
sorted_eigen_vectors[26][11] = 64'b1011111110111100100100110001001011001000101001011000001000110101;
sorted_eigen_vectors[26][12] = 64'b1011111110000110100110010010000110110010001100011010000010011100;
sorted_eigen_vectors[26][13] = 64'b0011111101101111000011110100101110101111111011100111000101101010;
sorted_eigen_vectors[26][14] = 64'b0011111101100101100001000110010001001111001010011011010110000000;
sorted_eigen_vectors[26][15] = 64'b0011111110001001010000100101001100011011000010110010000000100011;
sorted_eigen_vectors[26][16] = 64'b1011111111011011100000101100001101110100110010101000001001001101;
sorted_eigen_vectors[26][17] = 64'b1011111111001111000101101110100101011010010100111100101100111110;
sorted_eigen_vectors[26][18] = 64'b0011111111000000110101110011100010101100101011110101100010100000;
sorted_eigen_vectors[26][19] = 64'b1011111110111010000010110110010011000010001100001100111111001110;
sorted_eigen_vectors[26][20] = 64'b1011111101111111001111011011001011110111101011000010100011100100;
sorted_eigen_vectors[26][21] = 64'b1011111111011110011110000100111110010010111010000111110100111101;
sorted_eigen_vectors[26][22] = 64'b1011111111010100011100001001100111101001111011011110001100011110;
sorted_eigen_vectors[26][23] = 64'b1011111101111001001010101000100000010110001110110011100010001100;
sorted_eigen_vectors[26][24] = 64'b1011111110010010000101010110111010001001110011001001101101010110;
sorted_eigen_vectors[26][25] = 64'b1011111110010110010101101110000110011110110100100011101011010110;
sorted_eigen_vectors[26][26] = 64'b1011111110100111101100111101100111000000111001100101100101100000;
sorted_eigen_vectors[26][27] = 64'b1011111110011010001010010010110011110110011101011111001110000111;
sorted_eigen_vectors[26][28] = 64'b0011111110110111010001011101010000111011011000000001001100011100;
sorted_eigen_vectors[26][29] = 64'b0011111101111001111000111010101101100110111000100101001000001011;
sorted_eigen_vectors[26][30] = 64'b1011111101111000111011000011100100110101010110110110011000101100;
sorted_eigen_vectors[26][31] = 64'b0011111100111101011100101000011110001011100101010111101000010010;
sorted_eigen_vectors[27][0] = 64'b1011111111001110010011100000001101100111111010000101010011111011;
sorted_eigen_vectors[27][1] = 64'b1011111110011010001101111001010111000110011101011100101011010001;
sorted_eigen_vectors[27][2] = 64'b0011111101110111110010001011001010000101101000110000000001110101;
sorted_eigen_vectors[27][3] = 64'b0011111110101111110010111010001001100100011001111011011110011010;
sorted_eigen_vectors[27][4] = 64'b1011111110110011100110110110000111100110100110010000001000000111;
sorted_eigen_vectors[27][5] = 64'b0011111110100000011010111011100111000001111101011111110101101000;
sorted_eigen_vectors[27][6] = 64'b0011111110110100000011010111100000101011001000010100110100110001;
sorted_eigen_vectors[27][7] = 64'b0011111111000110110011101101111010000100001001101011100000110111;
sorted_eigen_vectors[27][8] = 64'b0011111110111111101101011101001011101000110111111000011010101101;
sorted_eigen_vectors[27][9] = 64'b0011111110110100000110010110001110100100011100011001111101110011;
sorted_eigen_vectors[27][10] = 64'b1011111110100100110110110010000100010011111101000101111110001111;
sorted_eigen_vectors[27][11] = 64'b1011111111011101101111111001000110110011101000101000010000111100;
sorted_eigen_vectors[27][12] = 64'b1011111110100100011000110000000000100110000110100001100011011011;
sorted_eigen_vectors[27][13] = 64'b0011111111010010101100110101010000111101110001001011100111101001;
sorted_eigen_vectors[27][14] = 64'b1011111111000111000001001111100111011001101001100111111001111011;
sorted_eigen_vectors[27][15] = 64'b1011111110101010111110010000011110111001110100011000111111000100;
sorted_eigen_vectors[27][16] = 64'b0011111111011010110010101011101100011110101011100010010011000100;
sorted_eigen_vectors[27][17] = 64'b0011111111010010111010111101001101110011010101101001101010011001;
sorted_eigen_vectors[27][18] = 64'b1011111111010101011001001001111111111110111110111111111011110011;
sorted_eigen_vectors[27][19] = 64'b0011111111000010011100001001001010101000110011000010010100000110;
sorted_eigen_vectors[27][20] = 64'b1011111111001111000010100000111110111111110101100110110000001011;
sorted_eigen_vectors[27][21] = 64'b1011111111010001001110111010001011111100010001100011000101110110;
sorted_eigen_vectors[27][22] = 64'b0011111110000001101011101011000110010110010011110110010010011001;
sorted_eigen_vectors[27][23] = 64'b0011111101111000110110111010111010101101010001111110001110100001;
sorted_eigen_vectors[27][24] = 64'b0011111110010010000000110111010110001000101000101111100100011101;
sorted_eigen_vectors[27][25] = 64'b0011111110110010100011001101011100100010011110101001100000011000;
sorted_eigen_vectors[27][26] = 64'b1011111110010111011100110001000010110111001001111101000001000011;
sorted_eigen_vectors[27][27] = 64'b1011111110001000101010111100110110110000100000110110101001100101;
sorted_eigen_vectors[27][28] = 64'b1011111110010111010001001101001011011100100111111101000101101010;
sorted_eigen_vectors[27][29] = 64'b0011111101011111000111111000011011110000000110011001110010000100;
sorted_eigen_vectors[27][30] = 64'b1011111101101001011111110110111001100010110000111100000100110111;
sorted_eigen_vectors[27][31] = 64'b1011111100110001001011100001000110011111110000010011001101011111;
sorted_eigen_vectors[28][0] = 64'b0011111101101011100101010111100101010011010101100101010001110101;
sorted_eigen_vectors[28][1] = 64'b1011111111000011001101110111100110000111000010101011001000001111;
sorted_eigen_vectors[28][2] = 64'b1011111110000001100010110110010000100101000000100110011010010101;
sorted_eigen_vectors[28][3] = 64'b0011111111010000001111111100111000101010011000100110001101010011;
sorted_eigen_vectors[28][4] = 64'b0011111111001101101001101011010101100001100110101111000110111011;
sorted_eigen_vectors[28][5] = 64'b0011111111000111100101001110000000010111011001000010011110111101;
sorted_eigen_vectors[28][6] = 64'b1011111110110000111100000010100010101010101110001010001110100011;
sorted_eigen_vectors[28][7] = 64'b1011111111001000000010001111011011101101101000001001110011100110;
sorted_eigen_vectors[28][8] = 64'b1011111111010100000100101000110100000011000100100110101100100010;
sorted_eigen_vectors[28][9] = 64'b0011111110101000101010000000101100001011100011000100101000110011;
sorted_eigen_vectors[28][10] = 64'b1011111110110011010011010010100111001100100101101111000111000010;
sorted_eigen_vectors[28][11] = 64'b1011111111010001100001111100000110100101011000001010000000001100;
sorted_eigen_vectors[28][12] = 64'b1011111111001010110111001101010000110110100110100110101111011001;
sorted_eigen_vectors[28][13] = 64'b1011111110011011011111010110001111011010000100111000010100001111;
sorted_eigen_vectors[28][14] = 64'b0011111111000001010010010111001101101101011011010010100100010101;
sorted_eigen_vectors[28][15] = 64'b0011111110110100111011100010010100011010100010100101101010010111;
sorted_eigen_vectors[28][16] = 64'b1011111111000001101000100000111100110000011000110110100101000010;
sorted_eigen_vectors[28][17] = 64'b1011111111010010101111110011011010101010100001011101110011100000;
sorted_eigen_vectors[28][18] = 64'b0011111110101001110010111001011001101000111010100010010100110000;
sorted_eigen_vectors[28][19] = 64'b0011111101110010100000100111010001111011100100010110011000111100;
sorted_eigen_vectors[28][20] = 64'b1011111111100100010100000110101100010011100011000000101101111111;
sorted_eigen_vectors[28][21] = 64'b0011111110111011000010011010010011101111110100101011101100000001;
sorted_eigen_vectors[28][22] = 64'b0011111110011100110111001001011101100111010100101000100111100001;
sorted_eigen_vectors[28][23] = 64'b1011111110010010110100110111110001011000100000010000100100110110;
sorted_eigen_vectors[28][24] = 64'b1011111110100011011100010010000011010101001010000101100100010001;
sorted_eigen_vectors[28][25] = 64'b1011111110011000110010001110110100001000000110101101110101110110;
sorted_eigen_vectors[28][26] = 64'b0011111110010000101100101101000110111110110101100100000111101010;
sorted_eigen_vectors[28][27] = 64'b1011111110110110001110001010010010110001111010000000101100001011;
sorted_eigen_vectors[28][28] = 64'b1011111110100111010001011101010000001100001110101110010101001000;
sorted_eigen_vectors[28][29] = 64'b1011111101110010001001000010010000011011111110000101001010111111;
sorted_eigen_vectors[28][30] = 64'b1011111101111111010000100010100011100000000001100011001100110110;
sorted_eigen_vectors[28][31] = 64'b1011111101000101101010100100011101001101101110101011110001001001;
sorted_eigen_vectors[29][0] = 64'b1011111101111011101100010101001101011001010000010101011110010010;
sorted_eigen_vectors[29][1] = 64'b1011111111000010000011011100110000001111100000101111101111000001;
sorted_eigen_vectors[29][2] = 64'b1011111110101000111111111011101100110011011011001000100101101010;
sorted_eigen_vectors[29][3] = 64'b0011111111010000111101001110010001001001010101000011111011011010;
sorted_eigen_vectors[29][4] = 64'b0011111111001101111011011111010101011010101011111111011000100011;
sorted_eigen_vectors[29][5] = 64'b0011111111001011000110010010101000001100111001101100111010001111;
sorted_eigen_vectors[29][6] = 64'b1011111110110110010000000001101011000010111010001100101011100001;
sorted_eigen_vectors[29][7] = 64'b1011111111001011000010110111101010011000110010100001000001000101;
sorted_eigen_vectors[29][8] = 64'b1011111111001111100101011001100000101011001011110110000000111101;
sorted_eigen_vectors[29][9] = 64'b0011111110000111011001010100011100000101010111111100110000001110;
sorted_eigen_vectors[29][10] = 64'b1011111110111100100101001100000101011101111000001111100100010101;
sorted_eigen_vectors[29][11] = 64'b1011111111010011100100000110111100001110100000111110001101000011;
sorted_eigen_vectors[29][12] = 64'b1011111110111010000001000011010010000101001000001000100111000111;
sorted_eigen_vectors[29][13] = 64'b0011111110101000110000110001101100110010100100100101011000111010;
sorted_eigen_vectors[29][14] = 64'b0011111110101101000110110111000010010011000001101000000000000101;
sorted_eigen_vectors[29][15] = 64'b0011111110010111011101101011010110111011000011110101001000000001;
sorted_eigen_vectors[29][16] = 64'b1011111111010010000010111110110100011011111001110100001100000101;
sorted_eigen_vectors[29][17] = 64'b0011111111000101101111001001001101110000010101010111010111100111;
sorted_eigen_vectors[29][18] = 64'b1011111111001000010101110000000010010100111000101110100111000110;
sorted_eigen_vectors[29][19] = 64'b0011111111000011010101011111110110100111100111001011101010110100;
sorted_eigen_vectors[29][20] = 64'b0011111111100011011001000001100110111100001101010110010111110000;
sorted_eigen_vectors[29][21] = 64'b1011111111000010101011001101001011011100100100010001000101101100;
sorted_eigen_vectors[29][22] = 64'b0011111110110101110000111001101110110101001011010110100111101110;
sorted_eigen_vectors[29][23] = 64'b0011111110100111000110101001011101110001001110111110011011100100;
sorted_eigen_vectors[29][24] = 64'b0011111110101000111000000111110011100110000000100010011000111111;
sorted_eigen_vectors[29][25] = 64'b1011111101010110101101100010001100100001011010010010100010110001;
sorted_eigen_vectors[29][26] = 64'b1011111110000100101011110101000111110001100001001110101001100110;
sorted_eigen_vectors[29][27] = 64'b0011111110110000110011001111101101100101001110000010110000111010;
sorted_eigen_vectors[29][28] = 64'b0011111110011000010101110001010011001100101110011010100001110000;
sorted_eigen_vectors[29][29] = 64'b1011111100111101110010010001101100110110110110111011010000001011;
sorted_eigen_vectors[29][30] = 64'b0011111101110010011001000100011111101000110110001011110110000110;
sorted_eigen_vectors[29][31] = 64'b1011111101011000111011100001101010001110000000000100101110010000;
sorted_eigen_vectors[30][0] = 64'b1011111111011101000011010110010000101000001100100011001101100100;
sorted_eigen_vectors[30][1] = 64'b0011111110100101101000010011110100000011011011011001110111010011;
sorted_eigen_vectors[30][2] = 64'b1011111101101111011110011110011000001001100110011000001001010101;
sorted_eigen_vectors[30][3] = 64'b1011111110110010000100000111110101010110010110001010111111000110;
sorted_eigen_vectors[30][4] = 64'b0011111110111100100000001011000000010111011101000100101100110010;
sorted_eigen_vectors[30][5] = 64'b1011111110011011011000010010011101000001111011010111011100111001;
sorted_eigen_vectors[30][6] = 64'b1011111110011011000111000011000001000101001001100111100110111100;
sorted_eigen_vectors[30][7] = 64'b1011111110011000101001011110101111101000101110111100110011010011;
sorted_eigen_vectors[30][8] = 64'b1011111110011000000101001001011110011101110101011100110011111000;
sorted_eigen_vectors[30][9] = 64'b0011111101101001011100110011001010001110000101010110011000100001;
sorted_eigen_vectors[30][10] = 64'b0011111110100101111111111000001111101011101000111001110010110100;
sorted_eigen_vectors[30][11] = 64'b0011111110101110001010000110001111111101100010011110101110000010;
sorted_eigen_vectors[30][12] = 64'b0011111101010010111000000000010100000001001001110010111110110000;
sorted_eigen_vectors[30][13] = 64'b1011111110101000001100111001101101111011100010010110010111111011;
sorted_eigen_vectors[30][14] = 64'b0011111110011101101110101011000001101101111100111011110001101101;
sorted_eigen_vectors[30][15] = 64'b0011111110010001111000000100110011001111001101111011101101101010;
sorted_eigen_vectors[30][16] = 64'b0011111110001001010011111111100110101010010110110000000011011000;
sorted_eigen_vectors[30][17] = 64'b1011111110010011111001110001110010110100011001110110110101110111;
sorted_eigen_vectors[30][18] = 64'b0011111110101011100000101011011001111101110011011110010100001100;
sorted_eigen_vectors[30][19] = 64'b1011111110101001101111010110100010010001100111110010111101011101;
sorted_eigen_vectors[30][20] = 64'b0011111110100010000110011010011011100000010011000011011100111110;
sorted_eigen_vectors[30][21] = 64'b1011111110101111011101010101110010101111110110001001111111011100;
sorted_eigen_vectors[30][22] = 64'b0011111110111110101111100010101111101101010101110101111010011100;
sorted_eigen_vectors[30][23] = 64'b1011111110110100011010101101101101010011010000111000110011000101;
sorted_eigen_vectors[30][24] = 64'b0011111110110011001100110001110110010011000100000011000011111110;
sorted_eigen_vectors[30][25] = 64'b1011111111100001100010010001110110001110101001001001000001101111;
sorted_eigen_vectors[30][26] = 64'b1011111111100001001111100101101101100110000011000010110011111111;
sorted_eigen_vectors[30][27] = 64'b1011111110100011001010000101111101000101110010100111100011001101;
sorted_eigen_vectors[30][28] = 64'b1011111111010111010010000011000100110010110111111000011010001001;
sorted_eigen_vectors[30][29] = 64'b0011111101111000000110100101000000111100110111010000010111101101;
sorted_eigen_vectors[30][30] = 64'b1011111110100101000100001110011110010100100010000010111000110000;
sorted_eigen_vectors[30][31] = 64'b0011111101000110111010010001101110001110001101111110001101011010;
sorted_eigen_vectors[31][0] = 64'b1011111111011101011000101011100101001001101010111110100100110010;
sorted_eigen_vectors[31][1] = 64'b0011111110100111000010110100111111001000111010011100111110011000;
sorted_eigen_vectors[31][2] = 64'b1011111110000100110101001001011000111011000111100010010111010010;
sorted_eigen_vectors[31][3] = 64'b1011111110110000001101001011010100101101011101101101000111001010;
sorted_eigen_vectors[31][4] = 64'b0011111110111110011010010110001111011000001000001010011111111001;
sorted_eigen_vectors[31][5] = 64'b1011111110011101011010111011111010010001101100010010010100110110;
sorted_eigen_vectors[31][6] = 64'b1011111110011100011110001011001010100101011011001111111010011001;
sorted_eigen_vectors[31][7] = 64'b1011111110100010111100001010000110011000010110101011010110111001;
sorted_eigen_vectors[31][8] = 64'b1011111110010101100111001111011110000110000100011101110001001010;
sorted_eigen_vectors[31][9] = 64'b1011111101110111101011000100101100011101011001000011110011001010;
sorted_eigen_vectors[31][10] = 64'b0011111110010101111000010110011111011010100001100000111110100110;
sorted_eigen_vectors[31][11] = 64'b0011111110101001010010011101001001011100110100010100000010000101;
sorted_eigen_vectors[31][12] = 64'b0011111110001100101010111100110010001100100110001010000001100000;
sorted_eigen_vectors[31][13] = 64'b1011111110001000011001101100011100110011111100010010111010011111;
sorted_eigen_vectors[31][14] = 64'b0011111110011100101101011111011001001001100011010110100011010011;
sorted_eigen_vectors[31][15] = 64'b0011111110001100011100010110000100001011110001001101001100111100;
sorted_eigen_vectors[31][16] = 64'b0011111110000101100101110110110000001010011111110110010011011000;
sorted_eigen_vectors[31][17] = 64'b0011111100011111100110101101110000101001011111001111000010011111;
sorted_eigen_vectors[31][18] = 64'b1011111101111101100001110001010110101100011101110001010100101100;
sorted_eigen_vectors[31][19] = 64'b1011111101010011001010000110110110011101101111110011010111011000;
sorted_eigen_vectors[31][20] = 64'b1011111110010101011011110011110101001001010001011100101001011101;
sorted_eigen_vectors[31][21] = 64'b0011111110000100101001000101001111011010001001000101101010111000;
sorted_eigen_vectors[31][22] = 64'b0011111110001010001000101000111000111000101001001011111101110111;
sorted_eigen_vectors[31][23] = 64'b1011111110010100011001011001000100110001001010110010111111001001;
sorted_eigen_vectors[31][24] = 64'b0011111110011001010010100111000000101010011100100111010011111100;
sorted_eigen_vectors[31][25] = 64'b1011111111011100011011011100111110000111100000110101001110101001;
sorted_eigen_vectors[31][26] = 64'b0011111111100010001100001101011101011001100110110100010010010111;
sorted_eigen_vectors[31][27] = 64'b0011111111000000011000000010111001101001101010010100011111100110;
sorted_eigen_vectors[31][28] = 64'b0011111111011110001001000000110111001110110000011101111011101011;
sorted_eigen_vectors[31][29] = 64'b1011111110010111001011100001101001011110011011100011010100111011;
sorted_eigen_vectors[31][30] = 64'b0011111110010000100000010001001010010101000100000000010010000010;
sorted_eigen_vectors[31][31] = 64'b1011111100110100011110111101111100101100000011010111011101101111;      
    end
endmodule
