//`timescale 1ns / 1ps
//       file_sample_input = $fopen("train_sample.txt", "r");
//       if (file_sample_input == 0) begin
//       $display("FILE IS NULL");
//       $finish;
      // end
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.05.2024 09:28:12
// Design Name: 
// Module Name: nsl_ids_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module nsl_ids_tb;
//Parameters
    parameter PC_NUM = 32, MAJ_PC_NUM = 10,MIN_PC_NUM = 5, FP_SIZE = 64;
        
        // Inputs and Outputs
   logic clk, reset;
    real sorted_eigen_values [0:PC_NUM -1];
    real sorted_eigen_vectors [0:PC_NUM-1][0:PC_NUM-1];
    real input_samples [0:PC_NUM -1];
    real ids_out;
    //logic ids_out_f;
    
    //Instatiating the DUT
    nsl_ids #(.PC_NUM(PC_NUM), .MAJ_PC_NUM(MAJ_PC_NUM), .MIN_PC_NUM(MIN_PC_NUM), .FP_SIZE(FP_SIZE))
    dut(
      //  .clk(clk), .reset(reset),
        .sorted_eigen_values(sorted_eigen_values),   // Defining an array made up of (PC_NUM) elements each of (FP_SIZE) bits
        .sorted_eigen_vectors(sorted_eigen_vectors), // Defining an array made up of (PC_NUM * PC_NUM) elements each of (FP_SIZE) bits
        .input_samples(input_samples),               // Defining an array made up of (PC_NUM) elements each of (FP_SIZE) bits 
        .ids_out(ids_out)
    );
    
//    // Read data from CSV file and apply it to inputs
//   initial begin
   
//       // Variables for reading CSV file
//       integer file_eigen_values;
//       integer file_eigen_vectors;
//       integer file_sample_input;
       
//       bit [FP_SIZE-1:0] eigen_value_dec;
//       bit [FP_SIZE-1:0] eigen_vector_dec;
//       bit [FP_SIZE-1:0] sample_input_dec;

//       // Open the CSV files for reading 
//       file_eigen_values = $fopen("\Post PCA inputs\sorted_eig_val", "r");
//       file_eigen_vectors = $fopen("\Post PCA inputs\sorted_eig_vec", "r");
//       file_sample_input = $fopen("\Post PCA inputs\train_sample", "r");
       
//       // Read input samples
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           $fscanf(file_sample_input, "%d,", sample_input_dec);
//           input_samples[i] = $bitstoreal(sample_input_dec);
//       end
       
//       // Read sorted eigen values
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           $fscanf(file_eigen_values, "%d,", eigen_value_dec);
//           sorted_eigen_values[i] = $bitstoreal(eigen_value_dec);
//       end

//       // Read sorted eigen vectors
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           for (int j = 0; j < PC_NUM; j = j + 1) begin
//               $fscanf(file_eigen_vectors, "%d,", eigen_vector_dec);
//               sorted_eigen_vectors[i][j] = $bitstoreal(eigen_vector_dec);
//           end
//       end

//       // Close the CSV files
//       $fclose(file_eigen_values);
//       $fclose(file_eigen_vectors);
//       $fclose(file_sample_input);
       
//timeunit 1ns;

//timeprecision 100ps;
       
       // Read eigen_values  data from file
   initial begin
   
//---------------------------------------------- CLOCK ASSERTIONS ----------------------------------------------------------
$display($time, " << Starting the Simulation >>");
    reset = 1'b1;
    clk = 1'b1;

    #50 reset = ~reset; 
//       integer file_sample_input;
//       integer file_eigen_values;
//       integer file_eigen_vectors;
       
//       real sample_input_dec;
//       real sorted_eigen_value_dec;
//       real sorted_eigen_vector_dec;
       
//       file_sample_input = $fopen("train_sample.csv", "r");
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           $fscanf(file_sample_input, "%d,", sample_input_dec);
//           input_samples[i] = $realtobits(sample_input_dec);
//       end
//       $fclose(file_sample_input); 
         

//       file_eigen_values = $fopen("sorted_eig_val.csv", "r");
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           $fscanf(file_eigen_values, "%d\n", sorted_eigen_value_dec);
//           sorted_eigen_values[i] = $realtobits(sorted_eigen_value_dec);
//       end
//       $fclose(file_eigen_values);

//       // Read long_vector data from file
//       file_eigen_vectors = $fopen("sorted_eig_vec.csv", "r");
//       for (int i = 0; i < PC_NUM; i = i + 1) begin
//           for (int j = 0; j < PC_NUM; j = j + 1) begin
//               $fscanf(file_eigen_vectors, "%d,", sorted_eigen_vector_dec);
//               sorted_eigen_vectors[i][j] = $realtobits(sorted_eigen_vector_dec);
//           end
//           // Skip the newline character at the end of each line
//           $fgetc(file_eigen_vectors);
//       end
//       $fclose(file_eigen_vectors);
      
      // Manually input values for input_samples
//    input_samples[0] = 64'b;
//    input_samples[1] = 64'b;
//--------------------------------- ATTACK SAMPLE FOR TESTING ---------------------------------------------------------------------------
//input_samples[0] = -0.129;
//input_samples[1] = -0.0314;
//input_samples[2] = -0.0661;
//input_samples[3] = -0.008620000000000001;
//input_samples[4] = -0.0999;
//input_samples[5] = -0.0279;
//input_samples[6] = -0.0155;
//input_samples[7] = -0.0451;
//input_samples[8] = -0.0333;
//input_samples[9] = -0.0169;
//input_samples[10] = -0.0342;
//input_samples[11] = -0.0236;
//input_samples[12] = -0.0555;
//input_samples[13] = 1.86;
//input_samples[14] = -0.36;
//input_samples[15] = 10.5;
//input_samples[16] = 11.4;
//input_samples[17] = -0.218;
//input_samples[18] = -0.221;
//input_samples[19] = -6.37;
//input_samples[20] = 0.28300000000000003;
//input_samples[21] = -0.465;
//input_samples[22] = 1.06;
//input_samples[23] = -1.77;
//input_samples[24] = -2.2;
//input_samples[25] = 0.0768;
//input_samples[26] = -0.479;
//input_samples[27] = -0.37799999999999995;
//input_samples[28] = 10.7;
//input_samples[29] = 17.5;
//input_samples[30] = -0.239;
//input_samples[31] = -0.233;

//--------------------------------- NORMAL SAMPLE FOR TESTTING ---------------------------------------------------------------------------
input_samples[0] = 0.0;
input_samples[1] = 0.0;
input_samples[2] = 1.0;
input_samples[3] = 0.0;
input_samples[4] = 0.0;
input_samples[5] = 0.0;
input_samples[6] = 0.0;
input_samples[7] = 0.0;
input_samples[8] = 0.0;
input_samples[9] = 0.0;
input_samples[10] = 0.0;
input_samples[11] = 0.0;
input_samples[12] = 0.0;
input_samples[13] = 0.0;
input_samples[14] = 0.0;
input_samples[15] = 0.0;
input_samples[16] = 0.0;
input_samples[17] = 0.88;
input_samples[18] = 0.0;
input_samples[19] = 0.0;
input_samples[20] = 0.0;
input_samples[21] = 0.0;
input_samples[22] = 0.0;
input_samples[23] = 0.0;
input_samples[24] = 0.0;
input_samples[25] = 0.6;
input_samples[26] = 2.0;
input_samples[27] = 0.0;
input_samples[28] = 0.0;
input_samples[29] = 0.0;
input_samples[30] = 0.0;
input_samples[31] = 0.0;


// Manually input values for sorted_eigen_values
sorted_eigen_values[0] = 4.007806153051598;
sorted_eigen_values[1] = 3.4662555042130507;
sorted_eigen_values[2] = 2.8590554335101905;
sorted_eigen_values[3] = 2.165422469619612;
sorted_eigen_values[4] = 1.9519983988087384;
sorted_eigen_values[5] = 1.5178085791262554;
sorted_eigen_values[6] = 1.3806933792110334;
sorted_eigen_values[7] = 1.34498213436319;
sorted_eigen_values[8] = 1.2491960719323412;
sorted_eigen_values[9] = 1.1341483545317097;
sorted_eigen_values[10] = 1.07607103592575;
sorted_eigen_values[11] = 1.043396333266135;
sorted_eigen_values[12] = 0.9978889787474562;
sorted_eigen_values[13] = 0.9897702736466968;
sorted_eigen_values[14] = 0.913647561839854;
sorted_eigen_values[15] = 0.8586762570609626;
sorted_eigen_values[16] = 0.7304777916681624;
sorted_eigen_values[17] = 0.6379129459010248;
sorted_eigen_values[18] = 0.5856154479707647;
sorted_eigen_values[19] = 0.5528774723065824;
sorted_eigen_values[20] = 0.5404923008142296;
sorted_eigen_values[21] = 0.4878278385496541;
sorted_eigen_values[22] = 0.39812281826152296;
sorted_eigen_values[23] = 0.2666997035609402;
sorted_eigen_values[24] = 0.24062141130919126;
sorted_eigen_values[25] = 0.1872934136948884;
sorted_eigen_values[26] = 0.1211492172159305;
sorted_eigen_values[27] = 0.11538843979272374;
sorted_eigen_values[28] = 0.10728430560602754;
sorted_eigen_values[29] = 0.0551239435206308;
sorted_eigen_values[30] = 0.016239457836917482;
sorted_eigen_values[31] = 0.0005317594984161127;

    // Repeat for all PC_NUM elements

// Manually input values for sorted_eigen_vectors
sorted_eigen_vectors[0][0] = -0.02702249373494993;
sorted_eigen_vectors[0][1] = -0.27812949583950225;
sorted_eigen_vectors[0][2] = -0.044430671901207516;
sorted_eigen_vectors[0][3] = -0.11001503564049171;
sorted_eigen_vectors[0][4] = 0.08373350413901327;
sorted_eigen_vectors[0][5] = 0.28962240778723125;
sorted_eigen_vectors[0][6] = 0.13121840789974742;
sorted_eigen_vectors[0][7] = 0.004792633705085637;
sorted_eigen_vectors[0][8] = 0.048119643538991605;
sorted_eigen_vectors[0][9] = -0.20457565982504752;
sorted_eigen_vectors[0][10] = -0.21829374810735327;
sorted_eigen_vectors[0][11] = 0.3241412087497341;
sorted_eigen_vectors[0][12] = 0.14772751398594502;
sorted_eigen_vectors[0][13] = 0.021991088103831206;
sorted_eigen_vectors[0][14] = 0.014656921393525995;
sorted_eigen_vectors[0][15] = -0.021145395218187226;
sorted_eigen_vectors[0][16] = -0.11030885849412062;
sorted_eigen_vectors[0][17] = 0.24196879956840145;
sorted_eigen_vectors[0][18] = -0.3884178085896777;
sorted_eigen_vectors[0][19] = 0.28087113819172915;
sorted_eigen_vectors[0][20] = -0.14920112493903406;
sorted_eigen_vectors[0][21] = 0.34500363945591683;
sorted_eigen_vectors[0][22] = -0.3355166597141456;
sorted_eigen_vectors[0][23] = 0.09947358434628754;
sorted_eigen_vectors[0][24] = -0.013445588476697247;
sorted_eigen_vectors[0][25] = -0.09308989512151597;
sorted_eigen_vectors[0][26] = -0.0579229054325029;
sorted_eigen_vectors[0][27] = -0.012372714575816766;
sorted_eigen_vectors[0][28] = -0.05691199777683044;
sorted_eigen_vectors[0][29] = 7.549764112710317e-05;
sorted_eigen_vectors[0][30] = 0.004922393618113742;
sorted_eigen_vectors[0][31] = 0.0007862639347934516;
sorted_eigen_vectors[1][0] = 0.0026269784586696356;
sorted_eigen_vectors[1][1] = -0.03367287501411907;
sorted_eigen_vectors[1][2] = -0.007037381449339847;
sorted_eigen_vectors[1][3] = 0.019387463130287524;
sorted_eigen_vectors[1][4] = -0.0004521050609124148;
sorted_eigen_vectors[1][5] = 0.13925021231731552;
sorted_eigen_vectors[1][6] = -0.6236900018038957;
sorted_eigen_vectors[1][7] = 0.2448750225637377;
sorted_eigen_vectors[1][8] = 0.1418046318899627;
sorted_eigen_vectors[1][9] = -0.16402337408264656;
sorted_eigen_vectors[1][10] = 0.04731093589452867;
sorted_eigen_vectors[1][11] = 0.04951869900900829;
sorted_eigen_vectors[1][12] = 0.023202768164828295;
sorted_eigen_vectors[1][13] = -0.013319352092342777;
sorted_eigen_vectors[1][14] = -0.07708038417502677;
sorted_eigen_vectors[1][15] = 0.058240722360333674;
sorted_eigen_vectors[1][16] = 0.16039284938196002;
sorted_eigen_vectors[1][17] = -0.4245691241233319;
sorted_eigen_vectors[1][18] = -0.017102983302665756;
sorted_eigen_vectors[1][19] = 0.5015715434607814;
sorted_eigen_vectors[1][20] = 0.07966772985411923;
sorted_eigen_vectors[1][21] = -0.047459590382765454;
sorted_eigen_vectors[1][22] = 0.04109958812707805;
sorted_eigen_vectors[1][23] = 0.008409780165564342;
sorted_eigen_vectors[1][24] = 0.010423991845572644;
sorted_eigen_vectors[1][25] = -0.001399505361390401;
sorted_eigen_vectors[1][26] = 0.000715980567645858;
sorted_eigen_vectors[1][27] = 0.001505592977205236;
sorted_eigen_vectors[1][28] = -0.0037439386022227556;
sorted_eigen_vectors[1][29] = -0.0002710101310663373;
sorted_eigen_vectors[1][30] = -0.0001722683943087726;
sorted_eigen_vectors[1][31] = 0.00034362047076801533;
sorted_eigen_vectors[2][0] = 0.002067818691324879;
sorted_eigen_vectors[2][1] = -0.06850927578448027;
sorted_eigen_vectors[2][2] = -0.10460214235292313;
sorted_eigen_vectors[2][3] = 0.055605665650372796;
sorted_eigen_vectors[2][4] = 0.01477165132337316;
sorted_eigen_vectors[2][5] = 0.14459401129210928;
sorted_eigen_vectors[2][6] = -0.6281533921324812;
sorted_eigen_vectors[2][7] = 0.18463602105096366;
sorted_eigen_vectors[2][8] = 0.10762314257976788;
sorted_eigen_vectors[2][9] = -0.0716995954673666;
sorted_eigen_vectors[2][10] = -0.01607042728530603;
sorted_eigen_vectors[2][11] = 0.006093640387732372;
sorted_eigen_vectors[2][12] = 0.01259827455088087;
sorted_eigen_vectors[2][13] = 0.012482674773353613;
sorted_eigen_vectors[2][14] = -0.008162744603771822;
sorted_eigen_vectors[2][15] = -0.029535244249531536;
sorted_eigen_vectors[2][16] = -0.1594135354553871;
sorted_eigen_vectors[2][17] = 0.3973364316268703;
sorted_eigen_vectors[2][18] = -0.013521963691952943;
sorted_eigen_vectors[2][19] = -0.5598361781408884;
sorted_eigen_vectors[2][20] = -0.12085426194757568;
sorted_eigen_vectors[2][21] = 0.0263527457030063;
sorted_eigen_vectors[2][22] = -0.021387338977708927;
sorted_eigen_vectors[2][23] = -0.01957683984359322;
sorted_eigen_vectors[2][24] = -0.006284760220143668;
sorted_eigen_vectors[2][25] = 0.009772272319635166;
sorted_eigen_vectors[2][26] = 0.005329552091986661;
sorted_eigen_vectors[2][27] = -0.002772194426139944;
sorted_eigen_vectors[2][28] = 0.0011291604327996205;
sorted_eigen_vectors[2][29] = -0.0007429228818481175;
sorted_eigen_vectors[2][30] = 0.0003025679499807726;
sorted_eigen_vectors[2][31] = -0.001083182572726828;
sorted_eigen_vectors[3][0] = -0.002167485241867769;
sorted_eigen_vectors[3][1] = -0.03235197713540865;
sorted_eigen_vectors[3][2] = -0.055823601579964716;
sorted_eigen_vectors[3][3] = -0.008582109427083333;
sorted_eigen_vectors[3][4] = -0.009512556320932864;
sorted_eigen_vectors[3][5] = 0.047602332952146595;
sorted_eigen_vectors[3][6] = -0.0435156425054125;
sorted_eigen_vectors[3][7] = -0.06451687224848779;
sorted_eigen_vectors[3][8] = 0.2217056296603864;
sorted_eigen_vectors[3][9] = 0.6067110719418395;
sorted_eigen_vectors[3][10] = -0.215642900550432;
sorted_eigen_vectors[3][11] = 0.10348759073330605;
sorted_eigen_vectors[3][12] = 0.039964250144721485;
sorted_eigen_vectors[3][13] = -0.018379756079943056;
sorted_eigen_vectors[3][14] = -0.1542273898955097;
sorted_eigen_vectors[3][15] = 0.6827380822711877;
sorted_eigen_vectors[3][16] = -0.019886649468035006;
sorted_eigen_vectors[3][17] = -0.05672909682977247;
sorted_eigen_vectors[3][18] = -0.10592417800598734;
sorted_eigen_vectors[3][19] = -0.04624376211348371;
sorted_eigen_vectors[3][20] = 0.023887975462155604;
sorted_eigen_vectors[3][21] = 0.02356417859371965;
sorted_eigen_vectors[3][22] = 0.007588546195761451;
sorted_eigen_vectors[3][23] = 0.053286959264141516;
sorted_eigen_vectors[3][24] = -0.0019060463117986375;
sorted_eigen_vectors[3][25] = -0.004825636178545783;
sorted_eigen_vectors[3][26] = -0.0017555372660914307;
sorted_eigen_vectors[3][27] = -0.0002956680479548149;
sorted_eigen_vectors[3][28] = -0.0009633732424207447;
sorted_eigen_vectors[3][29] = -0.00030264097615287643;
sorted_eigen_vectors[3][30] = 0.0005335055116945844;
sorted_eigen_vectors[3][31] = -0.002039004700992699;
sorted_eigen_vectors[4][0] = 0.008953918257974258;
sorted_eigen_vectors[4][1] = -0.06554459565133522;
sorted_eigen_vectors[4][2] = 0.039386553576197116;
sorted_eigen_vectors[4][3] = 0.0003040877013351283;
sorted_eigen_vectors[4][4] = -0.027621442053776226;
sorted_eigen_vectors[4][5] = 0.06486272357346455;
sorted_eigen_vectors[4][6] = -0.014701218677951397;
sorted_eigen_vectors[4][7] = -0.025662770348880034;
sorted_eigen_vectors[4][8] = -0.15200002291670994;
sorted_eigen_vectors[4][9] = 0.2328238182054517;
sorted_eigen_vectors[4][10] = 0.6971938721365217;
sorted_eigen_vectors[4][11] = 0.1764736105305319;
sorted_eigen_vectors[4][12] = 0.20939053758569756;
sorted_eigen_vectors[4][13] = 0.33948186661463353;
sorted_eigen_vectors[4][14] = -0.21365978818320389;
sorted_eigen_vectors[4][15] = -0.04784251361346319;
sorted_eigen_vectors[4][16] = -0.34705145660145487;
sorted_eigen_vectors[4][17] = -0.017642635387365296;
sorted_eigen_vectors[4][18] = -0.16982727438479636;
sorted_eigen_vectors[4][19] = 0.07438539015735757;
sorted_eigen_vectors[4][20] = -0.1179029130125862;
sorted_eigen_vectors[4][21] = -0.12549197097864126;
sorted_eigen_vectors[4][22] = 0.03166640165505293;
sorted_eigen_vectors[4][23] = -0.005009993970240852;
sorted_eigen_vectors[4][24] = 0.02620772809480789;
sorted_eigen_vectors[4][25] = 0.009377069314629716;
sorted_eigen_vectors[4][26] = -0.0012169142846607517;
sorted_eigen_vectors[4][27] = -0.008723787512065;
sorted_eigen_vectors[4][28] = -0.0006697734758222033;
sorted_eigen_vectors[4][29] = -0.0012610280677217219;
sorted_eigen_vectors[4][30] = -0.000651855554411114;
sorted_eigen_vectors[4][31] = -0.0003520347310810604;
sorted_eigen_vectors[5][0] = -0.005525858645822891;
sorted_eigen_vectors[5][1] = -0.04693774409608019;
sorted_eigen_vectors[5][2] = -0.03534688772157832;
sorted_eigen_vectors[5][3] = 0.0038269110059594358;
sorted_eigen_vectors[5][4] = 0.010684837638402082;
sorted_eigen_vectors[5][5] = 0.08704314704368422;
sorted_eigen_vectors[5][6] = -0.1039873191691063;
sorted_eigen_vectors[5][7] = -0.07477456804724551;
sorted_eigen_vectors[5][8] = 0.15735030666305838;
sorted_eigen_vectors[5][9] = 0.6051404513300102;
sorted_eigen_vectors[5][10] = -0.22068225789519824;
sorted_eigen_vectors[5][11] = 0.1333072061107564;
sorted_eigen_vectors[5][12] = 0.001634093953437625;
sorted_eigen_vectors[5][13] = -0.060004291047950076;
sorted_eigen_vectors[5][14] = 0.14388222096114986;
sorted_eigen_vectors[5][15] = -0.685446555178378;
sorted_eigen_vectors[5][16] = 0.0018502178683417918;
sorted_eigen_vectors[5][17] = -0.10045724711101464;
sorted_eigen_vectors[5][18] = -0.03938350608844349;
sorted_eigen_vectors[5][19] = 0.04659085946912027;
sorted_eigen_vectors[5][20] = -0.010598854571223379;
sorted_eigen_vectors[5][21] = -0.06306251925162056;
sorted_eigen_vectors[5][22] = 0.019436524732652647;
sorted_eigen_vectors[5][23] = 0.04871580798397178;
sorted_eigen_vectors[5][24] = 0.005200572213717127;
sorted_eigen_vectors[5][25] = -0.010719202007929206;
sorted_eigen_vectors[5][26] = 0.002292706487299615;
sorted_eigen_vectors[5][27] = -0.0056046917270982;
sorted_eigen_vectors[5][28] = 0.0003478710104280906;
sorted_eigen_vectors[5][29] = 0.00023122681478255727;
sorted_eigen_vectors[5][30] = -0.0003960513365657888;
sorted_eigen_vectors[5][31] = -0.0017759972102174702;
sorted_eigen_vectors[6][0] = -0.0081491196189142;
sorted_eigen_vectors[6][1] = -0.17447188829716573;
sorted_eigen_vectors[6][2] = -0.4102665892315246;
sorted_eigen_vectors[6][3] = -0.09601566032340914;
sorted_eigen_vectors[6][4] = -0.08960129697184083;
sorted_eigen_vectors[6][5] = -0.23978992711311506;
sorted_eigen_vectors[6][6] = -0.01974943183239849;
sorted_eigen_vectors[6][7] = 0.25044077473440574;
sorted_eigen_vectors[6][8] = -0.37628000516209714;
sorted_eigen_vectors[6][9] = 0.08852932992740799;
sorted_eigen_vectors[6][10] = -0.10795998650131604;
sorted_eigen_vectors[6][11] = 0.024163590327659842;
sorted_eigen_vectors[6][12] = 0.048718619936911504;
sorted_eigen_vectors[6][13] = 0.020358009268331652;
sorted_eigen_vectors[6][14] = -0.009703995909207591;
sorted_eigen_vectors[6][15] = 0.006039064175968405;
sorted_eigen_vectors[6][16] = -0.0005028765143426599;
sorted_eigen_vectors[6][17] = 0.012634726903057256;
sorted_eigen_vectors[6][18] = 0.03912206101348005;
sorted_eigen_vectors[6][19] = 0.053244102969305644;
sorted_eigen_vectors[6][20] = 0.004894239473669784;
sorted_eigen_vectors[6][21] = -0.01424882787345829;
sorted_eigen_vectors[6][22] = 0.01056519288951662;
sorted_eigen_vectors[6][23] = 0.039103529104827964;
sorted_eigen_vectors[6][24] = -0.0004327692976503548;
sorted_eigen_vectors[6][25] = -0.001885219655660864;
sorted_eigen_vectors[6][26] = 0.00027630110457597956;
sorted_eigen_vectors[6][27] = -8.283416139526509e-05;
sorted_eigen_vectors[6][28] = 0.0005905780000549367;
sorted_eigen_vectors[6][29] = 0.00040179649043673143;
sorted_eigen_vectors[6][30] = -0.0014299937744925214;
sorted_eigen_vectors[6][31] = 0.7016665190057249;
sorted_eigen_vectors[7][0] = -0.011280218871434992;
sorted_eigen_vectors[7][1] = -0.17225888158182764;
sorted_eigen_vectors[7][2] = -0.3435001606978468;
sorted_eigen_vectors[7][3] = -0.024735980238699887;
sorted_eigen_vectors[7][4] = -0.01640567017723505;
sorted_eigen_vectors[7][5] = 0.06043122675621749;
sorted_eigen_vectors[7][6] = 0.0402513796465375;
sorted_eigen_vectors[7][7] = -0.20001928222355161;
sorted_eigen_vectors[7][8] = 0.3600597004224544;
sorted_eigen_vectors[7][9] = -0.05184856131109487;
sorted_eigen_vectors[7][10] = 0.18187044295496135;
sorted_eigen_vectors[7][11] = -0.10510439739488961;
sorted_eigen_vectors[7][12] = -0.05343079252024041;
sorted_eigen_vectors[7][13] = -0.03928187689705196;
sorted_eigen_vectors[7][14] = 0.029187753919371368;
sorted_eigen_vectors[7][15] = 0.022464892399130968;
sorted_eigen_vectors[7][16] = -0.08252553066235607;
sorted_eigen_vectors[7][17] = 0.2364839166835299;
sorted_eigen_vectors[7][18] = 0.4616157702246637;
sorted_eigen_vectors[7][19] = 0.22912943346511025;
sorted_eigen_vectors[7][20] = -0.10151833476276463;
sorted_eigen_vectors[7][21] = -0.07492349873386946;
sorted_eigen_vectors[7][22] = 0.08616036609455982;
sorted_eigen_vectors[7][23] = 0.5196590709935786;
sorted_eigen_vectors[7][24] = -0.01645448703555549;
sorted_eigen_vectors[7][25] = -0.042475283107461535;
sorted_eigen_vectors[7][26] = -0.005832407413002639;
sorted_eigen_vectors[7][27] = -0.0027081235564310434;
sorted_eigen_vectors[7][28] = 0.00031568798558642106;
sorted_eigen_vectors[7][29] = -0.0022071316290225955;
sorted_eigen_vectors[7][30] = -0.00028942368827680553;
sorted_eigen_vectors[7][31] = 0.0015440017438448294;
sorted_eigen_vectors[8][0] = -0.012656872081340174;
sorted_eigen_vectors[8][1] = -0.21290058999916345;
sorted_eigen_vectors[8][2] = -0.4049063401758341;
sorted_eigen_vectors[8][3] = -0.03308439782938224;
sorted_eigen_vectors[8][4] = -0.009592917355657057;
sorted_eigen_vectors[8][5] = 0.03972972632736708;
sorted_eigen_vectors[8][6] = 0.058318146927982685;
sorted_eigen_vectors[8][7] = -0.1831898462045448;
sorted_eigen_vectors[8][8] = 0.3028564825008108;
sorted_eigen_vectors[8][9] = -0.022484113848555642;
sorted_eigen_vectors[8][10] = 0.13170238248938204;
sorted_eigen_vectors[8][11] = -0.05788100409950735;
sorted_eigen_vectors[8][12] = -0.08977820743522429;
sorted_eigen_vectors[8][13] = -0.0436836550583951;
sorted_eigen_vectors[8][14] = 0.036705801348135454;
sorted_eigen_vectors[8][15] = -0.00024365917425321631;
sorted_eigen_vectors[8][16] = -0.027301828487680913;
sorted_eigen_vectors[8][17] = 0.015737141689334395;
sorted_eigen_vectors[8][18] = 0.053380413364800816;
sorted_eigen_vectors[8][19] = 0.08113891047999432;
sorted_eigen_vectors[8][20] = 0.014740611692001469;
sorted_eigen_vectors[8][21] = 0.009875233652674014;
sorted_eigen_vectors[8][22] = -0.0587190364457124;
sorted_eigen_vectors[8][23] = -0.7780301366461254;
sorted_eigen_vectors[8][24] = 0.030355680477714232;
sorted_eigen_vectors[8][25] = 0.07190269377556327;
sorted_eigen_vectors[8][26] = 0.022307829552189358;
sorted_eigen_vectors[8][27] = 0.012235318086374597;
sorted_eigen_vectors[8][28] = 0.00851922008257379;
sorted_eigen_vectors[8][29] = 0.0033250943885130588;
sorted_eigen_vectors[8][30] = -0.0037550390571881053;
sorted_eigen_vectors[8][31] = 0.015624958165160888;
sorted_eigen_vectors[9][0] = -0.008416613327086124;
sorted_eigen_vectors[9][1] = -0.18000643960524232;
sorted_eigen_vectors[9][2] = -0.4197140604983773;
sorted_eigen_vectors[9][3] = -0.09756008334198847;
sorted_eigen_vectors[9][4] = -0.09021398322032083;
sorted_eigen_vectors[9][5] = -0.23563418005451756;
sorted_eigen_vectors[9][6] = -0.014865582652868047;
sorted_eigen_vectors[9][7] = 0.2403884833651897;
sorted_eigen_vectors[9][8] = -0.3600196313693195;
sorted_eigen_vectors[9][9] = 0.07979522606253758;
sorted_eigen_vectors[9][10] = -0.09879041104394186;
sorted_eigen_vectors[9][11] = 0.021503038491343003;
sorted_eigen_vectors[9][12] = 0.044189260641384;
sorted_eigen_vectors[9][13] = 0.01829734926504199;
sorted_eigen_vectors[9][14] = -0.008436360446797799;
sorted_eigen_vectors[9][15] = 0.00474920627654392;
sorted_eigen_vectors[9][16] = 0.002455426346610426;
sorted_eigen_vectors[9][17] = 0.0036901895168354204;
sorted_eigen_vectors[9][18] = 0.0321989337372028;
sorted_eigen_vectors[9][19] = 0.047437714469213646;
sorted_eigen_vectors[9][20] = 0.0068982657916355685;
sorted_eigen_vectors[9][21] = -0.013030346096797919;
sorted_eigen_vectors[9][22] = 0.008826048717655636;
sorted_eigen_vectors[9][23] = 0.027961073734073773;
sorted_eigen_vectors[9][24] = -0.0008650471852292774;
sorted_eigen_vectors[9][25] = -0.0016292911803775824;
sorted_eigen_vectors[9][26] = -0.0017283183783753427;
sorted_eigen_vectors[9][27] = -0.0003800686754575456;
sorted_eigen_vectors[9][28] = 0.00206296262913272;
sorted_eigen_vectors[9][29] = 4.193165201937982e-06;
sorted_eigen_vectors[9][30] = 0.0009701064504095145;
sorted_eigen_vectors[9][31] = -0.712179197277211;
sorted_eigen_vectors[10][0] = -0.004296433149463887;
sorted_eigen_vectors[10][1] = -0.09301256507333547;
sorted_eigen_vectors[10][2] = -0.04474477082029684;
sorted_eigen_vectors[10][3] = 0.050913921518722115;
sorted_eigen_vectors[10][4] = 0.10193356782415068;
sorted_eigen_vectors[10][5] = 0.29224907916493303;
sorted_eigen_vectors[10][6] = 0.043983108583960095;
sorted_eigen_vectors[10][7] = -0.2322366362643446;
sorted_eigen_vectors[10][8] = -0.12968269228003906;
sorted_eigen_vectors[10][9] = -0.132242406032523;
sorted_eigen_vectors[10][10] = -0.3126880690289034;
sorted_eigen_vectors[10][11] = 0.17907636280481828;
sorted_eigen_vectors[10][12] = 0.37890114338842246;
sorted_eigen_vectors[10][13] = 0.3399392458601293;
sorted_eigen_vectors[10][14] = -0.4137477771522329;
sorted_eigen_vectors[10][15] = -0.06430143217066453;
sorted_eigen_vectors[10][16] = 0.20201192797249054;
sorted_eigen_vectors[10][17] = -0.0908048673316289;
sorted_eigen_vectors[10][18] = 0.3490200139360532;
sorted_eigen_vectors[10][19] = -0.1353114459265384;
sorted_eigen_vectors[10][20] = 0.010088976601083842;
sorted_eigen_vectors[10][21] = -0.16068724167872067;
sorted_eigen_vectors[10][22] = 0.112944836282478;
sorted_eigen_vectors[10][23] = -0.08217273503951812;
sorted_eigen_vectors[10][24] = 0.0027216333512583885;
sorted_eigen_vectors[10][25] = 0.03785709358454;
sorted_eigen_vectors[10][26] = 0.0162092425486823;
sorted_eigen_vectors[10][27] = 0.002609551723871808;
sorted_eigen_vectors[10][28] = 0.012130017787365721;
sorted_eigen_vectors[10][29] = 0.0007432473266666597;
sorted_eigen_vectors[10][30] = -0.001749197223063407;
sorted_eigen_vectors[10][31] = -0.0016145711861073077;
sorted_eigen_vectors[11][0] = 0.0017648688769941558;
sorted_eigen_vectors[11][1] = -0.01985709812672651;
sorted_eigen_vectors[11][2] = 0.0070020672905648255;
sorted_eigen_vectors[11][3] = 0.0015223055131738732;
sorted_eigen_vectors[11][4] = 0.004031467506438393;
sorted_eigen_vectors[11][5] = 0.024961701329063644;
sorted_eigen_vectors[11][6] = 0.0024798897294898937;
sorted_eigen_vectors[11][7] = -0.023604484734772373;
sorted_eigen_vectors[11][8] = -0.014190497891196422;
sorted_eigen_vectors[11][9] = 0.029517442821726525;
sorted_eigen_vectors[11][10] = 0.08111190575746002;
sorted_eigen_vectors[11][11] = -0.3590152826080505;
sorted_eigen_vectors[11][12] = 0.7391866546544947;
sorted_eigen_vectors[11][13] = -0.5539427258525809;
sorted_eigen_vectors[11][14] = -0.02151485717053503;
sorted_eigen_vectors[11][15] = -0.017051180537957032;
sorted_eigen_vectors[11][16] = -0.014081643736748481;
sorted_eigen_vectors[11][17] = -0.005329983420547162;
sorted_eigen_vectors[11][18] = -0.06729683767821172;
sorted_eigen_vectors[11][19] = 0.003206993976280403;
sorted_eigen_vectors[11][20] = -0.049383236660592765;
sorted_eigen_vectors[11][21] = 0.007459269909217584;
sorted_eigen_vectors[11][22] = 0.012125596714057118;
sorted_eigen_vectors[11][23] = -0.017763172579623437;
sorted_eigen_vectors[11][24] = -0.003416758063994449;
sorted_eigen_vectors[11][25] = 0.0043993589725318215;
sorted_eigen_vectors[11][26] = 0.005559170978844449;
sorted_eigen_vectors[11][27] = -0.0014923145515788685;
sorted_eigen_vectors[11][28] = -0.0038470852188498446;
sorted_eigen_vectors[11][29] = 6.447908984075955e-05;
sorted_eigen_vectors[11][30] = 2.1044021193742525e-05;
sorted_eigen_vectors[11][31] = -5.894592357666707e-05;
sorted_eigen_vectors[12][0] = -0.005088620998649089;
sorted_eigen_vectors[12][1] = -0.17177172792444342;
sorted_eigen_vectors[12][2] = -0.3376878035158214;
sorted_eigen_vectors[12][3] = -0.05102339450290672;
sorted_eigen_vectors[12][4] = -0.034697895880189414;
sorted_eigen_vectors[12][5] = 0.040389576872789115;
sorted_eigen_vectors[12][6] = 0.09508019362128162;
sorted_eigen_vectors[12][7] = -0.1821499857103335;
sorted_eigen_vectors[12][8] = 0.16524088116581337;
sorted_eigen_vectors[12][9] = -0.19605511053316377;
sorted_eigen_vectors[12][10] = 0.11675888722002012;
sorted_eigen_vectors[12][11] = -0.019877679720214675;
sorted_eigen_vectors[12][12] = -0.058088922744738015;
sorted_eigen_vectors[12][13] = -0.012005175854831471;
sorted_eigen_vectors[12][14] = -0.02775281856716034;
sorted_eigen_vectors[12][15] = -0.05199449731657581;
sorted_eigen_vectors[12][16] = 0.1498459375110705;
sorted_eigen_vectors[12][17] = -0.4654961341181418;
sorted_eigen_vectors[12][18] = -0.4554401616512733;
sorted_eigen_vectors[12][19] = -0.4227152495346553;
sorted_eigen_vectors[12][20] = 0.1049631012901573;
sorted_eigen_vectors[12][21] = -0.04506239231250773;
sorted_eigen_vectors[12][22] = 0.07020531577421298;
sorted_eigen_vectors[12][23] = 0.27967805896595904;
sorted_eigen_vectors[12][24] = -0.009090551730828771;
sorted_eigen_vectors[12][25] = -0.010641729521007448;
sorted_eigen_vectors[12][26] = -0.0045694294008726925;
sorted_eigen_vectors[12][27] = -0.007639251671446047;
sorted_eigen_vectors[12][28] = 0.008272958437177859;
sorted_eigen_vectors[12][29] = -0.0029020214143907776;
sorted_eigen_vectors[12][30] = 0.0043252786464244766;
sorted_eigen_vectors[12][31] = 0.013944922672763937;
sorted_eigen_vectors[13][0] = 0.12930633737682126;
sorted_eigen_vectors[13][1] = 0.16130050712702643;
sorted_eigen_vectors[13][2] = -0.09076605579209047;
sorted_eigen_vectors[13][3] = -0.2990483711369147;
sorted_eigen_vectors[13][4] = 0.4966976719796876;
sorted_eigen_vectors[13][5] = 0.01593815855649134;
sorted_eigen_vectors[13][6] = 0.03977168312804918;
sorted_eigen_vectors[13][7] = 0.14204652908167326;
sorted_eigen_vectors[13][8] = 0.04653253211581921;
sorted_eigen_vectors[13][9] = 0.04900392280281063;
sorted_eigen_vectors[13][10] = 0.03602848439655803;
sorted_eigen_vectors[13][11] = -0.1339013633880835;
sorted_eigen_vectors[13][12] = -0.06726003144792396;
sorted_eigen_vectors[13][13] = 0.0057452152363081715;
sorted_eigen_vectors[13][14] = -0.21393079081908697;
sorted_eigen_vectors[13][15] = -0.060192778619213225;
sorted_eigen_vectors[13][16] = -0.018392524783189552;
sorted_eigen_vectors[13][17] = -0.013804218745129479;
sorted_eigen_vectors[13][18] = 0.006105827149093985;
sorted_eigen_vectors[13][19] = -0.01056392531556755;
sorted_eigen_vectors[13][20] = 0.007557513765853131;
sorted_eigen_vectors[13][21] = 0.14473186495193746;
sorted_eigen_vectors[13][22] = 0.03314023456209582;
sorted_eigen_vectors[13][23] = 0.013972824447738754;
sorted_eigen_vectors[13][24] = 0.07856589731239831;
sorted_eigen_vectors[13][25] = 0.005577151719735081;
sorted_eigen_vectors[13][26] = -0.005249857943834541;
sorted_eigen_vectors[13][27] = 0.024333916795615407;
sorted_eigen_vectors[13][28] = 0.019362866444246788;
sorted_eigen_vectors[13][29] = 0.6932337398772357;
sorted_eigen_vectors[13][30] = 0.04882865332895342;
sorted_eigen_vectors[13][31] = -4.1059123798355676e-05;
sorted_eigen_vectors[14][0] = 0.13685285986456797;
sorted_eigen_vectors[14][1] = 0.18026668924144928;
sorted_eigen_vectors[14][2] = -0.10152677425077007;
sorted_eigen_vectors[14][3] = -0.296245767506754;
sorted_eigen_vectors[14][4] = 0.4836557423364156;
sorted_eigen_vectors[14][5] = 0.0328131759271938;
sorted_eigen_vectors[14][6] = 0.045930709094100214;
sorted_eigen_vectors[14][7] = 0.14735320728416607;
sorted_eigen_vectors[14][8] = 0.045195454044017785;
sorted_eigen_vectors[14][9] = 0.045623809955549884;
sorted_eigen_vectors[14][10] = 0.033354753380326126;
sorted_eigen_vectors[14][11] = -0.12024822354868263;
sorted_eigen_vectors[14][12] = -0.06468462721209958;
sorted_eigen_vectors[14][13] = 0.00041087585595755803;
sorted_eigen_vectors[14][14] = -0.20301865567313296;
sorted_eigen_vectors[14][15] = -0.05714347607416074;
sorted_eigen_vectors[14][16] = -0.02035612803770944;
sorted_eigen_vectors[14][17] = -0.0012526188339400765;
sorted_eigen_vectors[14][18] = -0.003610990708526482;
sorted_eigen_vectors[14][19] = -0.002419758921405245;
sorted_eigen_vectors[14][20] = 0.02009098169674683;
sorted_eigen_vectors[14][21] = 0.11019407126581145;
sorted_eigen_vectors[14][22] = 0.04451184846364404;
sorted_eigen_vectors[14][23] = -0.001125099627289311;
sorted_eigen_vectors[14][24] = -0.08369564129896896;
sorted_eigen_vectors[14][25] = 0.0023904012986586697;
sorted_eigen_vectors[14][26] = -0.008792442264088499;
sorted_eigen_vectors[14][27] = -0.04241883228129952;
sorted_eigen_vectors[14][28] = -0.007894291287890522;
sorted_eigen_vectors[14][29] = -0.7051147303607354;
sorted_eigen_vectors[14][30] = -0.049203123388969074;
sorted_eigen_vectors[14][31] = 0.0002500572993668624;
sorted_eigen_vectors[15][0] = -0.004436082160828022;
sorted_eigen_vectors[15][1] = -0.0809600888538704;
sorted_eigen_vectors[15][2] = -0.034890294255225954;
sorted_eigen_vectors[15][3] = 0.4921196985605779;
sorted_eigen_vectors[15][4] = 0.3109791045838071;
sorted_eigen_vectors[15][5] = -0.25226346340194405;
sorted_eigen_vectors[15][6] = 0.07993141582902343;
sorted_eigen_vectors[15][7] = 0.15149331092974247;
sorted_eigen_vectors[15][8] = 0.1323964939930784;
sorted_eigen_vectors[15][9] = -0.0107795755747889;
sorted_eigen_vectors[15][10] = 0.04186996345079795;
sorted_eigen_vectors[15][11] = 0.16335917388831037;
sorted_eigen_vectors[15][12] = 0.06287791914995419;
sorted_eigen_vectors[15][13] = -0.029692304120092182;
sorted_eigen_vectors[15][14] = -0.03347040032414197;
sorted_eigen_vectors[15][15] = -0.015826703250062246;
sorted_eigen_vectors[15][16] = 0.06310443539922897;
sorted_eigen_vectors[15][17] = -0.019854200441710483;
sorted_eigen_vectors[15][18] = 0.0030002018405940684;
sorted_eigen_vectors[15][19] = -0.019587420143635965;
sorted_eigen_vectors[15][20] = -0.07994314519747907;
sorted_eigen_vectors[15][21] = 0.023755434503397614;
sorted_eigen_vectors[15][22] = -0.03623424478946652;
sorted_eigen_vectors[15][23] = 0.027238125071388574;
sorted_eigen_vectors[15][24] = 0.10192815583854983;
sorted_eigen_vectors[15][25] = 0.0854677340047767;
sorted_eigen_vectors[15][26] = -0.18228568259935674;
sorted_eigen_vectors[15][27] = 0.6563169193936436;
sorted_eigen_vectors[15][28] = 0.0877535029580827;
sorted_eigen_vectors[15][29] = -0.05358845243031962;
sorted_eigen_vectors[15][30] = 0.045018156132307856;
sorted_eigen_vectors[15][31] = 6.388852436716092e-05;
sorted_eigen_vectors[16][0] = -0.012909523304185865;
sorted_eigen_vectors[16][1] = -0.07200092427668163;
sorted_eigen_vectors[16][2] = -0.043178964221557536;
sorted_eigen_vectors[16][3] = 0.4928666564589183;
sorted_eigen_vectors[16][4] = 0.30232742100642906;
sorted_eigen_vectors[16][5] = -0.24094852144234266;
sorted_eigen_vectors[16][6] = 0.08726196550333062;
sorted_eigen_vectors[16][7] = 0.1657578412710153;
sorted_eigen_vectors[16][8] = 0.145704998764843;
sorted_eigen_vectors[16][9] = -0.014786951655621081;
sorted_eigen_vectors[16][10] = 0.052631485664868416;
sorted_eigen_vectors[16][11] = 0.17457563295448966;
sorted_eigen_vectors[16][12] = 0.08048141970511091;
sorted_eigen_vectors[16][13] = -0.017600181894357924;
sorted_eigen_vectors[16][14] = -0.020281040080182704;
sorted_eigen_vectors[16][15] = -0.011885589617580062;
sorted_eigen_vectors[16][16] = 0.07401786688436922;
sorted_eigen_vectors[16][17] = 0.03901551686410069;
sorted_eigen_vectors[16][18] = -0.010687562891629138;
sorted_eigen_vectors[16][19] = -0.005468233980691224;
sorted_eigen_vectors[16][20] = 0.08287909884611094;
sorted_eigen_vectors[16][21] = -0.015232603055064315;
sorted_eigen_vectors[16][22] = -0.005422381926860297;
sorted_eigen_vectors[16][23] = -7.78832424929083e-05;
sorted_eigen_vectors[16][24] = -0.1257991226626349;
sorted_eigen_vectors[16][25] = -0.04974432193691782;
sorted_eigen_vectors[16][26] = 0.17051767775916424;
sorted_eigen_vectors[16][27] = -0.6547580128211569;
sorted_eigen_vectors[16][28] = -0.09078227732322484;
sorted_eigen_vectors[16][29] = 0.04910171853089972;
sorted_eigen_vectors[16][30] = -0.04766363597006282;
sorted_eigen_vectors[16][31] = -0.00031096229423297953;
sorted_eigen_vectors[17][0] = -0.4672908923507345;
sorted_eigen_vectors[17][1] = 0.04603396011459258;
sorted_eigen_vectors[17][2] = -0.007564045148290788;
sorted_eigen_vectors[17][3] = -0.08778960376447299;
sorted_eigen_vectors[17][4] = 0.1173014786215067;
sorted_eigen_vectors[17][5] = -0.01516199857752969;
sorted_eigen_vectors[17][6] = -0.03791164085121239;
sorted_eigen_vectors[17][7] = -0.05891425406809524;
sorted_eigen_vectors[17][8] = -0.04052977109055913;
sorted_eigen_vectors[17][9] = -0.004607519468528582;
sorted_eigen_vectors[17][10] = 0.02164709803027257;
sorted_eigen_vectors[17][11] = 0.07787432218188366;
sorted_eigen_vectors[17][12] = 0.003935325443562912;
sorted_eigen_vectors[17][13] = -0.048033327805566475;
sorted_eigen_vectors[17][14] = 0.054179250611946415;
sorted_eigen_vectors[17][15] = 0.016790405606893877;
sorted_eigen_vectors[17][16] = -0.036881473918418305;
sorted_eigen_vectors[17][17] = -0.02729043039015531;
sorted_eigen_vectors[17][18] = 0.03513823375931591;
sorted_eigen_vectors[17][19] = -0.0070280108199204695;
sorted_eigen_vectors[17][20] = 0.02498135500765529;
sorted_eigen_vectors[17][21] = 0.013592728470931945;
sorted_eigen_vectors[17][22] = -0.04658990881456385;
sorted_eigen_vectors[17][23] = 0.03784650976354707;
sorted_eigen_vectors[17][24] = -0.05938768401882642;
sorted_eigen_vectors[17][25] = 0.4513638646880177;
sorted_eigen_vectors[17][26] = -0.036396989844599645;
sorted_eigen_vectors[17][27] = -0.09209026769487624;
sorted_eigen_vectors[17][28] = -0.0490518470691733;
sorted_eigen_vectors[17][29] = -0.042402293767796986;
sorted_eigen_vectors[17][30] = 0.7141804640103834;
sorted_eigen_vectors[17][31] = 0.0009965027253868515;
sorted_eigen_vectors[18][0] = -0.4646012293156691;
sorted_eigen_vectors[18][1] = 0.044876307612361416;
sorted_eigen_vectors[18][2] = -0.007158662553028808;
sorted_eigen_vectors[18][3] = -0.09220283890053566;
sorted_eigen_vectors[18][4] = 0.11741074772752336;
sorted_eigen_vectors[18][5] = -0.015893723854584103;
sorted_eigen_vectors[18][6] = -0.04018552915874685;
sorted_eigen_vectors[18][7] = -0.0651133970440723;
sorted_eigen_vectors[18][8] = -0.04217156243908;
sorted_eigen_vectors[18][9] = -0.007365320765808948;
sorted_eigen_vectors[18][10] = 0.019768518267036093;
sorted_eigen_vectors[18][11] = 0.08251104270482285;
sorted_eigen_vectors[18][12] = 0.0043361601918071755;
sorted_eigen_vectors[18][13] = -0.04977917281474921;
sorted_eigen_vectors[18][14] = 0.053901819873501206;
sorted_eigen_vectors[18][15] = 0.016358682581581567;
sorted_eigen_vectors[18][16] = -0.0381485452002048;
sorted_eigen_vectors[18][17] = -0.027332306498975646;
sorted_eigen_vectors[18][18] = 0.025786534916595855;
sorted_eigen_vectors[18][19] = -0.005977405682947026;
sorted_eigen_vectors[18][20] = 0.02303884769436444;
sorted_eigen_vectors[18][21] = 0.026666923231772326;
sorted_eigen_vectors[18][22] = -0.05575349066469207;
sorted_eigen_vectors[18][23] = 0.05314087061716081;
sorted_eigen_vectors[18][24] = -0.0424701573829984;
sorted_eigen_vectors[18][25] = 0.4957994776856465;
sorted_eigen_vectors[18][26] = -0.008361852731991144;
sorted_eigen_vectors[18][27] = 0.008648079549431168;
sorted_eigen_vectors[18][28] = -0.015432653772308355;
sorted_eigen_vectors[18][29] = 0.048062015330835955;
sorted_eigen_vectors[18][30] = -0.6918035266459246;
sorted_eigen_vectors[18][31] = -0.0014815862268919393;
sorted_eigen_vectors[19][0] = -0.02844479331026724;
sorted_eigen_vectors[19][1] = 0.24667999526585596;
sorted_eigen_vectors[19][2] = -0.19546683463858694;
sorted_eigen_vectors[19][3] = 0.15944384423293356;
sorted_eigen_vectors[19][4] = -0.0759150653998839;
sorted_eigen_vectors[19][5] = 0.4533476868956817;
sorted_eigen_vectors[19][6] = 0.15641582392090275;
sorted_eigen_vectors[19][7] = 0.23502190355921304;
sorted_eigen_vectors[19][8] = -0.09210538429109816;
sorted_eigen_vectors[19][9] = 0.061403692201067124;
sorted_eigen_vectors[19][10] = 0.12715042800554602;
sorted_eigen_vectors[19][11] = 0.08556840755083574;
sorted_eigen_vectors[19][12] = -0.05313823490635504;
sorted_eigen_vectors[19][13] = -0.11369163040326755;
sorted_eigen_vectors[19][14] = 0.07386949481449474;
sorted_eigen_vectors[19][15] = 0.024005631811354684;
sorted_eigen_vectors[19][16] = 0.1030774450724011;
sorted_eigen_vectors[19][17] = 0.021301901830373123;
sorted_eigen_vectors[19][18] = 0.03267041667635062;
sorted_eigen_vectors[19][19] = -0.01743764871883804;
sorted_eigen_vectors[19][20] = 0.05339143856400276;
sorted_eigen_vectors[19][21] = -0.02565664723709488;
sorted_eigen_vectors[19][22] = 0.03519372565861186;
sorted_eigen_vectors[19][23] = -0.032668790142454815;
sorted_eigen_vectors[19][24] = -0.6894293612622575;
sorted_eigen_vectors[19][25] = -0.045328245982752285;
sorted_eigen_vectors[19][26] = -0.05939897754405753;
sorted_eigen_vectors[19][27] = 0.12955773047799055;
sorted_eigen_vectors[19][28] = 0.048721912235867686;
sorted_eigen_vectors[19][29] = 0.08872916088493164;
sorted_eigen_vectors[19][30] = 0.0018804075021382504;
sorted_eigen_vectors[19][31] = 0.0005605721006140185;
sorted_eigen_vectors[20][0] = 0.023296680251460408;
sorted_eigen_vectors[20][1] = -0.2398477792462633;
sorted_eigen_vectors[20][2] = 0.19221614256322705;
sorted_eigen_vectors[20][3] = -0.16160312060289575;
sorted_eigen_vectors[20][4] = 0.052155947337404585;
sorted_eigen_vectors[20][5] = -0.4511087432494486;
sorted_eigen_vectors[20][6] = -0.157705065004752;
sorted_eigen_vectors[20][7] = -0.234862542703417;
sorted_eigen_vectors[20][8] = 0.10255712835016392;
sorted_eigen_vectors[20][9] = -0.0628726343037052;
sorted_eigen_vectors[20][10] = -0.1306588601816581;
sorted_eigen_vectors[20][11] = -0.08907901909060174;
sorted_eigen_vectors[20][12] = 0.054427182325060074;
sorted_eigen_vectors[20][13] = 0.1336246503606978;
sorted_eigen_vectors[20][14] = -0.09827557965197357;
sorted_eigen_vectors[20][15] = -0.037449224491685584;
sorted_eigen_vectors[20][16] = -0.14343607168565678;
sorted_eigen_vectors[20][17] = 0.003908751698318472;
sorted_eigen_vectors[20][18] = -0.08386667314223843;
sorted_eigen_vectors[20][19] = 0.05522394346425084;
sorted_eigen_vectors[20][20] = -0.03213664553165198;
sorted_eigen_vectors[20][21] = -0.0004924879507616416;
sorted_eigen_vectors[20][22] = 0.10845385954001481;
sorted_eigen_vectors[20][23] = -0.034743259724261025;
sorted_eigen_vectors[20][24] = -0.6759721915759555;
sorted_eigen_vectors[20][25] = -0.05284260854228788;
sorted_eigen_vectors[20][26] = -0.05100039197527489;
sorted_eigen_vectors[20][27] = 0.10220519644691443;
sorted_eigen_vectors[20][28] = 0.0059520460339748124;
sorted_eigen_vectors[20][29] = 0.06137796553806471;
sorted_eigen_vectors[20][30] = 0.002375644911440169;
sorted_eigen_vectors[20][31] = 0.000262546233837342;
sorted_eigen_vectors[21][0] = -0.06804858503272164;
sorted_eigen_vectors[21][1] = 0.015009790137171563;
sorted_eigen_vectors[21][2] = 0.009250975898807908;
sorted_eigen_vectors[21][3] = 0.11543806386841443;
sorted_eigen_vectors[21][4] = -0.1740204283633179;
sorted_eigen_vectors[21][5] = -0.03154690363709711;
sorted_eigen_vectors[21][6] = -0.005890825721125436;
sorted_eigen_vectors[21][7] = -0.09477711827723093;
sorted_eigen_vectors[21][8] = -0.08820366643870693;
sorted_eigen_vectors[21][9] = -0.04188352356206948;
sorted_eigen_vectors[21][10] = -0.03412084468350759;
sorted_eigen_vectors[21][11] = 0.11277699827384398;
sorted_eigen_vectors[21][12] = -0.34304971986706234;
sorted_eigen_vectors[21][13] = -0.4886671834956812;
sorted_eigen_vectors[21][14] = -0.7095627820659803;
sorted_eigen_vectors[21][15] = -0.12074466125878447;
sorted_eigen_vectors[21][16] = -0.1230686120034225;
sorted_eigen_vectors[21][17] = 0.07249053445847026;
sorted_eigen_vectors[21][18] = -0.06838343505402653;
sorted_eigen_vectors[21][19] = 0.057965364411871334;
sorted_eigen_vectors[21][20] = -0.06577287694467017;
sorted_eigen_vectors[21][21] = -0.09538111536145265;
sorted_eigen_vectors[21][22] = -0.0318591274827871;
sorted_eigen_vectors[21][23] = 0.003382006068597124;
sorted_eigen_vectors[21][24] = 0.011456537770405185;
sorted_eigen_vectors[21][25] = -0.0016632625919491793;
sorted_eigen_vectors[21][26] = 0.009707161199504783;
sorted_eigen_vectors[21][27] = -0.01869852793225243;
sorted_eigen_vectors[21][28] = 0.004158426901939216;
sorted_eigen_vectors[21][29] = 0.000182686438807196;
sorted_eigen_vectors[21][30] = 0.000322896294754875;
sorted_eigen_vectors[21][31] = -0.00029262914477038294;
sorted_eigen_vectors[22][0] = 0.2054973643346205;
sorted_eigen_vectors[22][1] = -0.008357509486910261;
sorted_eigen_vectors[22][2] = 0.002877046069042528;
sorted_eigen_vectors[22][3] = -0.1888994306132261;
sorted_eigen_vectors[22][4] = 0.28674737357527263;
sorted_eigen_vectors[22][5] = -0.02698698446767794;
sorted_eigen_vectors[22][6] = -0.10740062481035939;
sorted_eigen_vectors[22][7] = -0.2209231908672719;
sorted_eigen_vectors[22][8] = -0.1658275199545796;
sorted_eigen_vectors[22][9] = -0.01935296613712841;
sorted_eigen_vectors[22][10] = 0.08282910457454146;
sorted_eigen_vectors[22][11] = 0.2751518423999047;
sorted_eigen_vectors[22][12] = -0.042933123784171204;
sorted_eigen_vectors[22][13] = -0.21911211175424686;
sorted_eigen_vectors[22][14] = 0.2083357312765699;
sorted_eigen_vectors[22][15] = 0.11145773372293433;
sorted_eigen_vectors[22][16] = 0.2706005375163584;
sorted_eigen_vectors[22][17] = 0.16047536002446386;
sorted_eigen_vectors[22][18] = -0.09769325087579506;
sorted_eigen_vectors[22][19] = 0.02980996627041471;
sorted_eigen_vectors[22][20] = -0.11417804958593053;
sorted_eigen_vectors[22][21] = -0.6223569507377884;
sorted_eigen_vectors[22][22] = -0.1980143531907875;
sorted_eigen_vectors[22][23] = -0.003945717273197985;
sorted_eigen_vectors[22][24] = -0.025684040461386705;
sorted_eigen_vectors[22][25] = -0.010210692417658493;
sorted_eigen_vectors[22][26] = 0.06879518933247042;
sorted_eigen_vectors[22][27] = 0.041065273220154366;
sorted_eigen_vectors[22][28] = -0.07784309413641739;
sorted_eigen_vectors[22][29] = 0.018550470625530575;
sorted_eigen_vectors[22][30] = 0.002448142180141671;
sorted_eigen_vectors[22][31] = -0.0007479718344251895;
sorted_eigen_vectors[23][0] = 0.051552331395803994;
sorted_eigen_vectors[23][1] = 0.40340196385469757;
sorted_eigen_vectors[23][2] = -0.20332575579766385;
sorted_eigen_vectors[23][3] = 0.04801580651789738;
sorted_eigen_vectors[23][4] = -0.0213095972235888;
sorted_eigen_vectors[23][5] = -0.08275369333258639;
sorted_eigen_vectors[23][6] = -0.01740822139357918;
sorted_eigen_vectors[23][7] = -0.09464270734194626;
sorted_eigen_vectors[23][8] = 0.06998819325463727;
sorted_eigen_vectors[23][9] = -0.13430088460636794;
sorted_eigen_vectors[23][10] = -0.19661515347301214;
sorted_eigen_vectors[23][11] = 0.10929782872070615;
sorted_eigen_vectors[23][12] = 0.09803091399003916;
sorted_eigen_vectors[23][13] = 0.04459691518967024;
sorted_eigen_vectors[23][14] = 0.08254924135113186;
sorted_eigen_vectors[23][15] = 0.017944785099403983;
sorted_eigen_vectors[23][16] = -0.2368533253972469;
sorted_eigen_vectors[23][17] = 0.03878416302053911;
sorted_eigen_vectors[23][18] = -0.19011556349493056;
sorted_eigen_vectors[23][19] = 0.1195762338453987;
sorted_eigen_vectors[23][20] = -0.18396728522157393;
sorted_eigen_vectors[23][21] = -0.17955171544552895;
sorted_eigen_vectors[23][22] = 0.24279644950764606;
sorted_eigen_vectors[23][23] = -0.027038222811317413;
sorted_eigen_vectors[23][24] = 0.06433927566465757;
sorted_eigen_vectors[23][25] = 0.04678975092509838;
sorted_eigen_vectors[23][26] = -0.3660614383647652;
sorted_eigen_vectors[23][27] = -0.18757536055754492;
sorted_eigen_vectors[23][28] = 0.5221895120117089;
sorted_eigen_vectors[23][29] = 0.008895775090546324;
sorted_eigen_vectors[23][30] = -0.006353903222693865;
sorted_eigen_vectors[23][31] = 0.00020400631358698799;
sorted_eigen_vectors[24][0] = -0.016289503020282883;
sorted_eigen_vectors[24][1] = 0.41324453088320295;
sorted_eigen_vectors[24][2] = -0.20842425605504003;
sorted_eigen_vectors[24][3] = 0.06908928025568126;
sorted_eigen_vectors[24][4] = -0.055762720492549836;
sorted_eigen_vectors[24][5] = -0.0696343481016284;
sorted_eigen_vectors[24][6] = 0.021054803921583046;
sorted_eigen_vectors[24][7] = -0.012884426727265818;
sorted_eigen_vectors[24][8] = 0.11366069011782147;
sorted_eigen_vectors[24][9] = -0.1185515074105174;
sorted_eigen_vectors[24][10] = -0.19901709919276883;
sorted_eigen_vectors[24][11] = 0.025507469232467554;
sorted_eigen_vectors[24][12] = 0.09747435824453601;
sorted_eigen_vectors[24][13] = 0.09664612465807618;
sorted_eigen_vectors[24][14] = 0.021679890386449904;
sorted_eigen_vectors[24][15] = -0.007733560718176947;
sorted_eigen_vectors[24][16] = -0.31046123542691273;
sorted_eigen_vectors[24][17] = -0.034461821536459596;
sorted_eigen_vectors[24][18] = -0.12958404817146577;
sorted_eigen_vectors[24][19] = 0.07691093458507142;
sorted_eigen_vectors[24][20] = -0.11011883658511949;
sorted_eigen_vectors[24][21] = -0.13866121720133678;
sorted_eigen_vectors[24][22] = 0.11201029983855668;
sorted_eigen_vectors[24][23] = -0.004572846817863995;
sorted_eigen_vectors[24][24] = 0.012379196653908608;
sorted_eigen_vectors[24][25] = -0.010667820925559672;
sorted_eigen_vectors[24][26] = 0.3987095191926637;
sorted_eigen_vectors[24][27] = 0.18251791870824197;
sorted_eigen_vectors[24][28] = -0.5732611725699078;
sorted_eigen_vectors[24][29] = 0.01217730019736948;
sorted_eigen_vectors[24][30] = 0.006963558227846671;
sorted_eigen_vectors[24][31] = -0.001727572876858795;
sorted_eigen_vectors[25][0] = 0.0012519462923298147;
sorted_eigen_vectors[25][1] = -0.3363436712559021;
sorted_eigen_vectors[25][2] = 0.1830916843325197;
sorted_eigen_vectors[25][3] = -0.1241406434168221;
sorted_eigen_vectors[25][4] = 0.043365756901375924;
sorted_eigen_vectors[25][5] = 0.1390400758896725;
sorted_eigen_vectors[25][6] = 0.14993076348953482;
sorted_eigen_vectors[25][7] = 0.23216492426983504;
sorted_eigen_vectors[25][8] = 0.0355330231748302;
sorted_eigen_vectors[25][9] = -0.05487940182984378;
sorted_eigen_vectors[25][10] = -0.029198484747059557;
sorted_eigen_vectors[25][11] = 0.1855225395000331;
sorted_eigen_vectors[25][12] = -0.05987048105418336;
sorted_eigen_vectors[25][13] = -0.1657898748754839;
sorted_eigen_vectors[25][14] = 0.09882458068527539;
sorted_eigen_vectors[25][15] = 0.038880855418204296;
sorted_eigen_vectors[25][16] = -0.031108485677827074;
sorted_eigen_vectors[25][17] = 0.09593121918385913;
sorted_eigen_vectors[25][18] = -0.08220373948616297;
sorted_eigen_vectors[25][19] = 0.01403233978392735;
sorted_eigen_vectors[25][20] = -0.0722308752858614;
sorted_eigen_vectors[25][21] = -0.07025717977404874;
sorted_eigen_vectors[25][22] = 0.771911705800084;
sorted_eigen_vectors[25][23] = -0.06311540730350859;
sorted_eigen_vectors[25][24] = 0.07029911465892137;
sorted_eigen_vectors[25][25] = 0.10919877023826664;
sorted_eigen_vectors[25][26] = 0.10709693880675217;
sorted_eigen_vectors[25][27] = 0.03044126496767307;
sorted_eigen_vectors[25][28] = -0.045534934775584776;
sorted_eigen_vectors[25][29] = 0.0001591787403627466;
sorted_eigen_vectors[25][30] = 0.002109175505534147;
sorted_eigen_vectors[25][31] = -0.0009645304121338643;
sorted_eigen_vectors[26][0] = -0.0684933405678625;
sorted_eigen_vectors[26][1] = -0.2151463040238767;
sorted_eigen_vectors[26][2] = 0.1439273698779929;
sorted_eigen_vectors[26][3] = -0.09828951848848365;
sorted_eigen_vectors[26][4] = 0.015255501649741593;
sorted_eigen_vectors[26][5] = 0.09613898070312411;
sorted_eigen_vectors[26][6] = 0.2127407755150423;
sorted_eigen_vectors[26][7] = 0.41101242713236313;
sorted_eigen_vectors[26][8] = 0.19169227661307453;
sorted_eigen_vectors[26][9] = -0.07002444689576709;
sorted_eigen_vectors[26][10] = -0.16870287431383152;
sorted_eigen_vectors[26][11] = -0.11161916159245139;
sorted_eigen_vectors[26][12] = -0.011034262896103812;
sorted_eigen_vectors[26][13] = 0.0037914732233287804;
sorted_eigen_vectors[26][14] = 0.0026266059078838278;
sorted_eigen_vectors[26][15] = 0.012333535445023415;
sorted_eigen_vectors[26][16] = -0.42985617070556686;
sorted_eigen_vectors[26][17] = -0.2428867045451514;
sorted_eigen_vectors[26][18] = 0.1315680354297841;
sorted_eigen_vectors[26][19] = -0.10173635235770392;
sorted_eigen_vectors[26][20] = -0.007627200214083117;
sorted_eigen_vectors[26][21] = -0.4760931906366358;
sorted_eigen_vectors[26][22] = -0.3193726334061909;
sorted_eigen_vectors[26][23] = -0.006144076909278107;
sorted_eigen_vectors[26][24] = -0.01765988079128119;
sorted_eigen_vectors[26][25] = -0.02181580097072352;
sorted_eigen_vectors[26][26] = -0.04629402618154432;
sorted_eigen_vectors[26][27] = -0.025547697584886755;
sorted_eigen_vectors[26][28] = 0.09090925645439224;
sorted_eigen_vectors[26][29] = 0.006320638216625439;
sorted_eigen_vectors[26][30] = -0.006084655256665832;
sorted_eigen_vectors[26][31] = 0.0004493313714045998;
sorted_eigen_vectors[27][0] = -0.2367557771073406;
sorted_eigen_vectors[27][1] = -0.025602665174526976;
sorted_eigen_vectors[27][2] = 0.0058066342846246795;
sorted_eigen_vectors[27][3] = 0.062100481754767865;
sorted_eigen_vectors[27][4] = -0.07658969764543865;
sorted_eigen_vectors[27][5] = 0.032071881224505834;
sorted_eigen_vectors[27][6] = 0.07833052685719079;
sorted_eigen_vectors[27][7] = 0.17818814709375072;
sorted_eigen_vectors[27][8] = 0.12386816201572046;
sorted_eigen_vectors[27][9] = 0.0785124088739602;
sorted_eigen_vectors[27][10] = -0.040734323202001765;
sorted_eigen_vectors[27][11] = -0.4648174528356924;
sorted_eigen_vectors[27][12] = -0.039817814494243556;
sorted_eigen_vectors[27][13] = 0.2921953776557574;
sorted_eigen_vectors[27][14] = -0.17983935477694846;
sorted_eigen_vectors[27][15] = -0.052681199486670084;
sorted_eigen_vectors[27][16] = 0.41862371441;
sorted_eigen_vectors[27][17] = 0.2956436754560997;
sorted_eigen_vectors[27][18] = -0.3342666616517668;
sorted_eigen_vectors[27][19] = 0.1440604519087076;
sorted_eigen_vectors[27][20] = -0.24249455325193056;
sorted_eigen_vectors[27][21] = -0.26926493297721465;
sorted_eigen_vectors[27][22] = 0.008633983039475534;
sorted_eigen_vectors[27][23] = 0.006068880397372662;
sorted_eigen_vectors[27][24] = 0.017591320480954235;
sorted_eigen_vectors[27][25] = 0.0724615534951173;
sorted_eigen_vectors[27][26] = -0.02289987676518047;
sorted_eigen_vectors[27][27] = -0.012046439122447692;
sorted_eigen_vectors[27][28] = -0.02272347899993702;
sorted_eigen_vectors[27][29] = 0.0018996064904060203;
sorted_eigen_vectors[27][30] = -0.0031125217411657425;
sorted_eigen_vectors[27][31] = -0.0002621453311391543;
sorted_eigen_vectors[28][0] = 0.0033671731604934477;
sorted_eigen_vectors[28][1] = -0.15013045400463954;
sorted_eigen_vectors[28][2] = -0.008566648845135286;
sorted_eigen_vectors[28][3] = 0.25389436854452646;
sorted_eigen_vectors[28][4] = 0.23165004030114555;
sorted_eigen_vectors[28][5] = 0.18423081533575028;
sorted_eigen_vectors[28][6] = -0.06616453330992882;
sorted_eigen_vectors[28][7] = -0.1877735767641077;
sorted_eigen_vectors[28][8] = -0.3136322526931271;
sorted_eigen_vectors[28][9] = 0.048157067451161245;
sorted_eigen_vectors[28][10] = -0.07539616818298271;
sorted_eigen_vectors[28][11] = -0.2739109148992617;
sorted_eigen_vectors[28][12] = -0.20986416498348495;
sorted_eigen_vectors[28][13] = -0.026845512566869678;
sorted_eigen_vectors[28][14] = 0.1350540432270654;
sorted_eigen_vectors[28][15] = 0.08175880334816052;
sorted_eigen_vectors[28][16] = -0.1377581583281629;
sorted_eigen_vectors[28][17] = -0.2929207482588492;
sorted_eigen_vectors[28][18] = 0.05038137465187232;
sorted_eigen_vectors[28][19] = 0.0045189428429580035;
sorted_eigen_vectors[28][20] = -0.6348166829851464;
sorted_eigen_vectors[28][21] = 0.10561591010148776;
sorted_eigen_vectors[28][22] = 0.02818523948793395;
sorted_eigen_vectors[28][23] = -0.018384879018648454;
sorted_eigen_vectors[28][24] = -0.037972475071159306;
sorted_eigen_vectors[28][25] = -0.024203971500097638;
sorted_eigen_vectors[28][26] = 0.016307141564142848;
sorted_eigen_vectors[28][27] = -0.08680180877130908;
sorted_eigen_vectors[28][28] = -0.045454622738768935;
sorted_eigen_vectors[28][29] = -0.004428998042858621;
sorted_eigen_vectors[28][30] = -0.007631454151476194;
sorted_eigen_vectors[28][31] = -0.0006611679231890512;
sorted_eigen_vectors[29][0] = -0.0067609077269334;
sorted_eigen_vectors[29][1] = -0.1410460544338701;
sorted_eigen_vectors[29][2] = -0.04882607462629347;
sorted_eigen_vectors[29][3] = 0.26494700585406655;
sorted_eigen_vectors[29][4] = 0.23382441452115285;
sorted_eigen_vectors[29][5] = 0.21170545225105683;
sorted_eigen_vectors[29][6] = -0.08691565760163257;
sorted_eigen_vectors[29][7] = -0.21128780804076733;
sorted_eigen_vectors[29][8] = -0.2467527590622484;
sorted_eigen_vectors[29][9] = 0.011423640109546464;
sorted_eigen_vectors[29][10] = -0.11164482633555325;
sorted_eigen_vectors[29][11] = -0.3056905404806011;
sorted_eigen_vectors[29][12] = -0.10162666559384724;
sorted_eigen_vectors[29][13] = 0.04836354248361059;
sorted_eigen_vectors[29][14] = 0.05684997362845937;
sorted_eigen_vectors[29][15] = 0.02291377977583587;
sorted_eigen_vectors[29][16] = -0.28197791790903215;
sorted_eigen_vectors[29][17] = 0.16981738076258;
sorted_eigen_vectors[29][18] = -0.1901550986274982;
sorted_eigen_vectors[29][19] = 0.15106173214140528;
sorted_eigen_vectors[29][20] = 0.6059693027447661;
sorted_eigen_vectors[29][21] = -0.1458991600976661;
sorted_eigen_vectors[29][22] = 0.0850159947707778;
sorted_eigen_vectors[29][23] = 0.04512475259066465;
sorted_eigen_vectors[29][24] = 0.048587706639477535;
sorted_eigen_vectors[29][25] = -0.0013861983367342953;
sorted_eigen_vectors[29][26] = -0.010100021536904437;
sorted_eigen_vectors[29][27] = 0.06562777730157245;
sorted_eigen_vectors[29][28] = 0.02376968860190981;
sorted_eigen_vectors[29][29] = -0.00045449175273298896;
sorted_eigen_vectors[29][30] = 0.004490166565616409;
sorted_eigen_vectors[29][31] = -0.0015216121028102968;
sorted_eigen_vectors[30][0] = -0.4539423363246924;
sorted_eigen_vectors[30][1] = 0.04224577586029068;
sorted_eigen_vectors[30][2] = -0.003842305461873511;
sorted_eigen_vectors[30][3] = -0.07056411130969228;
sorted_eigen_vectors[30][4] = 0.11133862087835379;
sorted_eigen_vectors[30][5] = -0.026737798117543597;
sorted_eigen_vectors[30][6] = -0.026474718304251733;
sorted_eigen_vectors[30][7] = -0.02407044036858681;
sorted_eigen_vectors[30][8] = -0.023516053207868176;
sorted_eigen_vectors[30][9] = 0.003106688251744997;
sorted_eigen_vectors[30][10] = 0.042965052141704346;
sorted_eigen_vectors[30][11] = 0.05890190572696154;
sorted_eigen_vectors[30][12] = 0.0011520432350264722;
sorted_eigen_vectors[30][13] = -0.04726873286262997;
sorted_eigen_vectors[30][14] = 0.02903247519583057;
sorted_eigen_vectors[30][15] = 0.01745719923740855;
sorted_eigen_vectors[30][16] = 0.012359571944557874;
sorted_eigen_vectors[30][17] = -0.019436310301768477;
sorted_eigen_vectors[30][18] = 0.053731634957282365;
sorted_eigen_vectors[30][19] = -0.0502731969605452;
sorted_eigen_vectors[30][20] = 0.035351958160488625;
sorted_eigen_vectors[30][21] = -0.06144227644500664;
sorted_eigen_vectors[30][22] = 0.12008928818192505;
sorted_eigen_vectors[30][23] = -0.07975550444421049;
sorted_eigen_vectors[30][24] = 0.07499871101771659;
sorted_eigen_vectors[30][25] = -0.5479877267830612;
sorted_eigen_vectors[30][26] = -0.5388619416347921;
sorted_eigen_vectors[30][27] = -0.03741739012660759;
sorted_eigen_vectors[30][28] = -0.3637812611396858;
sorted_eigen_vectors[30][29] = 0.0058844694411290645;
sorted_eigen_vectors[30][30] = -0.04114459694036687;
sorted_eigen_vectors[30][31] = 0.0006991753147636934;
sorted_eigen_vectors[31][0] = -0.45915062136159;
sorted_eigen_vectors[31][1] = 0.04500817611270164;
sorted_eigen_vectors[31][2] = -0.010171102217799186;
sorted_eigen_vectors[31][3] = -0.06330425605739902;
sorted_eigen_vectors[31][4] = 0.11879562403251487;
sorted_eigen_vectors[31][5] = -0.028731324808437732;
sorted_eigen_vectors[31][6] = -0.027804175707614044;
sorted_eigen_vectors[31][7] = -0.0369921205977834;
sorted_eigen_vectors[31][8] = -0.021106593664139955;
sorted_eigen_vectors[31][9] = -0.005779546181897641;
sorted_eigen_vectors[31][10] = 0.02136766692412064;
sorted_eigen_vectors[31][11] = 0.04939134009384907;
sorted_eigen_vectors[31][12] = 0.013999555626540592;
sorted_eigen_vectors[31][13] = -0.011914783737800248;
sorted_eigen_vectors[31][14] = 0.028037880172043846;
sorted_eigen_vectors[31][15] = 0.013888128444344273;
sorted_eigen_vectors[31][16] = 0.010542720861780472;
sorted_eigen_vectors[31][17] = 0.00012056320917691814;
sorted_eigen_vectors[31][18] = -0.007208904898509599;
sorted_eigen_vectors[31][19] = -0.0011693067999546305;
sorted_eigen_vectors[31][20] = -0.02093215713234496;
sorted_eigen_vectors[31][21] = 0.010079054922738848;
sorted_eigen_vectors[31][22] = 0.012761221984504561;
sorted_eigen_vectors[31][23] = -0.019918697954196127;
sorted_eigen_vectors[31][24] = 0.02469802149845622;
sorted_eigen_vectors[31][25] = -0.44420231088343565;
sorted_eigen_vectors[31][26] = 0.5684620618941549;
sorted_eigen_vectors[31][27] = 0.12793522032967458;
sorted_eigen_vectors[31][28] = 0.4709505576242765;
sorted_eigen_vectors[31][29] = -0.0226368065009883;
sorted_eigen_vectors[31][30] = 0.016117372844750573;
sorted_eigen_vectors[31][31] = -0.00031255911385651754;
    
    end
    
    always begin
        #50 clk = ~clk; // Toggle the clock every 5 time units
    end
endmodule
